
module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   N599, g1289, g1882, g312, g452, g11257, g123, g207, g713, g1153,
         g1744, g1558, g695, g461, g940, g976, g709, g8432, g1092, g1574,
         g1864, g369, g1580, g1736, g1424, g1737, g1672, g1077, g1231, g4,
         g1104, g1304, g7290, g243, g1499, g1444, g1543, g315, g1534, g622,
         g1927, g1660, g278, g1436, g718, g8433, g554, g496, g11333, g981,
         g829, g1095, g704, g1265, g7302, g1786, g682, g8429, g1296, g7292,
         g327, g1389, g1371, g1956, g1955, g1675, g354, g113, g639, g1684,
         g1639, g1791, g248, g1707, g1759, g351, g1604, g1098, g932, g1896,
         g8282, g736, g8435, g1019, g745, g1419, g32, g1086, g1486, g1730,
         g1504, g1470, g822, g1678, g174, g1766, g1801, g186, g959, g1407,
         g1868, g1718, g396, g11265, g1015, g1415, g1227, g1721, g284, g426,
         g11256, g219, g1360, g806, g1428, g1564, g1741, g225, g281, g1308,
         g611, g1217, g1589, g1466, g1571, g1861, g1448, g1133, g1333, g153,
         g962, g486, g11331, g471, g1397, g1950, g8288, g756, g755, g1101,
         g549, g105, g1669, g1531, g1458, g572, g1011, g1411, g1074, g444,
         g11259, g1474, g1080, g1713, g333, g269, g401, g11266, g1857, g9,
         g664, g965, g1400, g309, g814, g231, g557, g869, g875, g1383, g158,
         g627, g1023, g259, g1327, g654, g293, g1346, g1633, g1753, g1508,
         g1240, g7297, g538, g11326, g416, g11269, g542, g11325, g1681, g374,
         g563, g1914, g8284, g530, g11328, g575, g1936, g1317, g1356, g357,
         g386, g11263, g1601, g166, g501, g11334, g262, g1840, g318, g794,
         g302, g342, g1250, g7299, g1163, g1032, g1432, g1453, g363, g330,
         g1157, g928, g261, g516, g11337, g254, g861, g1627, g1292, g7293,
         g290, g1583, g466, g1561, g1546, g287, g560, g617, g336, g456, g305,
         g345, g8, g255, g1945, g1738, g1478, g1690, g1482, g1110, g296, g1663,
         g700, g8431, g1762, g360, g192, g1657, g722, g566, g1089, g1071, g986,
         g971, g143, g1814, g1212, g1918, g1822, g237, g746, g1462, g178, g366,
         g837, g599, g1854, g944, g1941, g8287, g170, g1520, g686, g953, g1958,
         g1765, g1733, g7303, g1610, g1796, g1324, g1540, g491, g11332, g213,
         g1781, g1900, g1245, g7298, g148, g833, g1923, g8285, g936, g1314,
         g849, g1336, g272, g1806, g826, g1887, g8281, g968, g1137, g1891,
         g1255, g7300, g257, g874, g591, g731, g636, g1218, g605, g182, g950,
         g1129, g857, g448, g11258, g1828, g1727, g1592, g1703, g1932, g8286,
         g1624, g440, g11260, g476, g11338, g119, g668, g139, g1149, g263,
         g818, g1747, g802, g275, g1524, g1577, g810, g391, g11264, g658,
         g1386, g253, g1125, g201, g1280, g7295, g1083, g650, g1636, g853,
         g421, g11270, g956, g378, g1756, g841, g1027, g1003, g1403, g1145,
         g1107, g1223, g406, g11267, g1811, g1654, g197, g1595, g1537, g727,
         g8434, g798, g481, g11324, g1330, g845, g1512, g1490, g1166, g348,
         g1260, g7301, g260, g131, g258, g521, g11330, g1318, g1872, g677,
         g1549, g947, g1834, g1598, g1121, g1321, g506, g11335, g546, g1909,
         g1552, g1687, g1586, g324, g1141, g1341, g1710, g135, g525, g11329,
         g1607, g321, g1275, g11443, g1615, g382, g266, g1284, g7294, g673,
         g8428, g162, g411, g11268, g431, g11262, g1905, g8283, g1515, g1630,
         g991, g1300, g7291, g339, g256, g1750, g1440, g1666, g1528, g1351,
         g127, g1618, g1235, g7296, g299, g435, g11261, g1555, g995, g1621,
         g643, g1494, g1567, g691, g8430, g534, g11327, g1776, g569, g1160, g1,
         g511, g11336, g1724, g12, g1878, g4500, g5529, g4338, g8147, g6551,
         g10865, g8054, g7709, g4940, g6481, g6529, g10707, g6949, g8940,
         g10855, g6920, g6907, g6155, g6638, g11647, g6910, g6828, g10800,
         g8019, g6821, g11478, g6516, g8244, g8631, g10793, g5910, g2478,
         g10726, g6824, g9961, g6759, g6502, g10797, g4471, g10780, g11625,
         g11372, g10771, g11293, g8173, g6533, g8245, g10767, g6000, g4490,
         g4903, g10720, g6934, g6123, g6838, g4905, g10798, g10785, g7204,
         g6830, g8944, g5543, g8921, g6096, g6942, g6733, g6823, g4890, g3381,
         g10863, g8039, g6526, g10664, g7189, g8923, g5173, g4264, g6755,
         g11514, g4506, g4465, g6902, g6015, g11340, g6542, g6507, g5556,
         g8505, g11641, g10765, g11305, g6126, g8060, g7191, g6469, g4498,
         g6627, g4893, g5194, g6901, g8043, g6929, g8049, g6786, g6234, g10864,
         g8984, g10862, g10721, g8051, g6541, g10773, g8193, g6523, g5404,
         g11393, g4334, g6908, g8768, g8885, g6333, g6045, g7590, g6468,
         g10782, g6672, g6840, g5914, g7705, g6038, g6471, g11303, g10663,
         g8920, g4283, g4484, g5396, g8045, g7843, g6932, g6537, g4902, g6080,
         g6059, g4089, g5126, g10866, g11603, g6332, g4231, g11488, g6955,
         g5918, g6894, g4076, g6534, g6928, g6926, g8055, g11291, g6833, g6918,
         g6915, g6911, g7441, g5996, g8047, g6653, g6832, g11481, g6478, g6897,
         g6042, g4342, g4330, g11609, g10859, g6054, g6508, g6531, g8050,
         g11376, g8559, g7032, g4293, g5390, g8767, g4480, g11483, g5392,
         g10776, g6513, g9272, g10898, g8052, g4325, g8766, g6205, g8820,
         g9124, g6839, g6522, g10936, g11320, g6841, g8769, g6224, g11349,
         g6470, g5755, g6515, g10791, g7632, g11485, g6331, g8053, g5763,
         g6480, g6795, g8194, g8938, g4238, g8775, g4891, g11290, g6501, g6334,
         g10719, g4274, g8765, g6916, g11308, g10784, g6820, g4340, g6922,
         g6747, g11391, g8649, g9555, g6071, g10858, g8926, g4239, g11602,
         g8041, g8922, g5536, g11605, g8048, g6528, g6524, g7219, g8046,
         g11482, g4477, g6923, g4255, g8937, g6538, g11306, g7183, g6895,
         g6179, g9721, g8776, g6827, g4309, g7244, g7586, g7930, g11300,
         g10718, g5445, g6088, g6679, g11636, g9266, g11608, g8059, g8771,
         g6035, g6198, g8973, g6834, g5148, g7134, g10795, g10770, g8773,
         g3462, g7143, g8939, g8772, g6093, g6500, g8777, g6244, g11640,
         g11487, g9110, g11380, g9269, g11314, g9150, g11298, g7202, g6819,
         g6243, g6514, g6983, g4473, g8040, g6900, g8042, g6546, g5770, g8889,
         g10711, g11312, g6479, g5849, g6656, g6906, g10717, g8770, g6392,
         g6621, g11610, g11604, g11486, g7581, g10799, g6439, g7133, g8044,
         g8254, g11607, g6193, g4904, g11292, g6822, g6912, g6898, g5421,
         g6924, g11310, g11294, g6026, g8024, g8945, g6525, g5083, g7541,
         g10860, g11579, g11639, g6826, g7626, g6829, g7660, g10722, g8887,
         g11484, g6002, g11606, g6757, g6216, g8941, g4892, g6930, g8250,
         g6049, g8943, g10861, g8779, g6180, g8774, g8260, g6099, g6831, g6068,
         g7137, g6545, g7257, g6909, g8384, g11392, g6506, g8883, g6728,
         g10724, g4556, DFF_121_n1, DFF_122_n1, DFF_126_n1, DFF_136_n1,
         DFF_157_n1, DFF_168_n1, DFF_194_n1, DFF_228_n1, g8271, DFF_242_n1,
         DFF_275_n1, DFF_311_n1, DFF_319_n1, DFF_330_n1, DFF_336_n1,
         DFF_350_n1, DFF_384_n1, DFF_385_n1, DFF_436_n1, DFF_441_n1,
         DFF_445_n1, DFF_452_n1, DFF_489_n1, n517, n518, n519, n520, n521,
         n522, n524, n526, n527, n528, n529, n530, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n542, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n583, n592, n594, n595,
         n596, n597, n598, n599, n600, n602, n603, n604, n605, n606, n607,
         n609, n610, n611, n612, n614, n616, n617, n619, n620, n621, n622,
         n623, n624, n625, n627, n629, n630, n631, n632, n633, n634, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n661, n662, n665,
         n667, n668, n674, n675, n685, n687, n711, n712, n713, n715, n717,
         n718, n719, n720, n721, n725, n744, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1459, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1583, n1585, n1586, n1587, n1588,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1727, n1729, n1731, n1733,
         n1735, n1737, n1739, n1741, n1743, n1745, n1747, n1749, n1751, n1753,
         n1755, n1757, n1759, n1761, n1763, n1765, n1767, n1769, n1771, n1773,
         n1775, n1777, n1779, n1781, n1783, n1785, n1787, n1789, n1791, n1793,
         n1795, n1797, n1799, n1801, n1803, n1805, n1807, n1809, n1811, n1813,
         n1815, n1817, n1819, n1821, n1823, n1825, n1827, n1829, n1831, n1833,
         n1835, n1837, g5105, n1839, g5101, n1841, n1843, n1845, n1847, n1849,
         n1851, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n3016, n3017, n3018, n3019,
         n3020, n3022, n3023, n3024, n3025, n3026, n3027, n3029, n3030, n3031,
         n3033, n3034, n3035, n3036, n3037, n3038, n3040, n3041, n3042, n3044,
         n3045, n3046, n3047, n3048, n3050, n3051, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3061, n3062, n3064, n3065;
  assign g8565 = g6949;
  assign g8561 = g6920;
  assign g9451 = g9961;
  assign g8564 = g6942;
  assign test_so10 = g8984;
  assign g8563 = g6932;
  assign g8566 = g6955;
  assign g8562 = g6926;
  assign g5816 = g8271;
  assign g11489 = 1'b0;
  assign g8062 = g5105;
  assign g8061 = g5101;

  LSDNENX1 U1550 ( .D(g10722), .ENB(n1887), .Q(g10461) );
  LSDNENX1 U1551 ( .D(g10664), .ENB(n1886), .Q(g10379) );
  SDFFX1 DFF_0_Q_reg ( .D(g4556), .SI(test_si1), .SE(test_se), .CLK(CK), .Q(
        g1289), .QN() );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(test_se), .CLK(CK), .Q(g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(test_se), .CLK(CK), .Q(g312), 
        .QN() );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(test_se), .CLK(CK), .Q(g452), 
        .QN() );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(test_se), .CLK(CK), .Q(g123), 
        .QN() );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(test_se), .CLK(CK), .Q(g207), 
        .QN() );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(test_se), .CLK(CK), .Q(g713), 
        .QN() );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(test_se), .CLK(CK), .Q(g1153), 
        .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(test_se), .CLK(CK), .Q(g1744), .QN() );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(test_se), .CLK(CK), .Q(
        g1558), .QN() );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(test_se), .CLK(CK), .Q(g695), .QN() );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(test_se), .CLK(CK), .Q(g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(test_se), .CLK(CK), .Q(g940), 
        .QN(n1712) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(test_se), .CLK(CK), .Q(g976), .QN() );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(test_se), .CLK(CK), .Q(g709), 
        .QN(n1719) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(test_se), .CLK(CK), .Q(g1092), .QN() );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(test_se), .CLK(CK), .Q(
        g1574), .QN() );
  SDFFX1 DFF_18_Q_reg ( .D(g6795), .SI(g1574), .SE(test_se), .CLK(CK), .Q(
        g1864), .QN() );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(test_se), .CLK(CK), .Q(
        g369), .QN() );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(test_se), .CLK(CK), .Q(g1580), .QN() );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(test_se), .CLK(CK), .Q(
        g1736), .QN() );
  SDFFX1 DFF_22_Q_reg ( .D(g10663), .SI(g1736), .SE(test_se), .CLK(CK), .Q(
        n1637), .QN() );
  SDFFX1 DFF_23_Q_reg ( .D(g10782), .SI(n1637), .SE(test_se), .CLK(CK), .Q(
        n3065), .QN(n1590) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(test_se), .CLK(CK), .Q(
        g1424), .QN() );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(test_se), .CLK(CK), .Q(
        g1737), .QN() );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(test_se), .CLK(CK), .Q(
        g1672), .QN() );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(test_se), .CLK(CK), .Q(
        g1077), .QN() );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(test_se), .CLK(CK), .Q(
        g1231), .QN() );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(test_se), .CLK(CK), .Q(g4), 
        .QN() );
  SDFFX1 DFF_30_Q_reg ( .D(g6728), .SI(g4), .SE(test_se), .CLK(CK), .Q(g4177), 
        .QN() );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(test_se), .CLK(CK), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(test_se), .CLK(CK), .Q(
        g1304), .QN() );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(test_se), .CLK(CK), .Q(g243), .QN() );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(test_se), .CLK(CK), .Q(g1499), .QN() );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(test_se), .CLK(CK), .Q(
        g1444), .QN() );
  SDFFX1 DFF_37_Q_reg ( .D(n524), .SI(g1444), .SE(test_se), .CLK(CK), .Q(n3064), .QN(n1868) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(test_se), .CLK(CK), .Q(
        g4180), .QN() );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(test_se), .CLK(CK), .Q(
        g1543), .QN() );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(test_se), .CLK(CK), .Q(g315), 
        .QN() );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(test_se), .CLK(CK), .Q(g1534), .QN(n1632) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(test_se), .CLK(CK), .Q(g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(test_se), .CLK(CK), .Q(g1927), .QN() );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(test_se), .CLK(CK), .Q(
        g1660), .QN() );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(test_se), .CLK(CK), .Q(g278), .QN() );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(test_se), .CLK(CK), .Q(g1436), .QN() );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(test_se), .CLK(CK), .Q(g718), .QN() );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(test_se), .CLK(CK), .Q(g8985), .QN(n1669) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(test_se), .CLK(CK), .Q(
        g554), .QN() );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(test_se), .CLK(CK), .Q(g496), .QN(n1689) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(test_se), .CLK(CK), .Q(g981), .QN(n1720) );
  SDFFX1 DFF_53_Q_reg ( .D(n616), .SI(g981), .SE(test_se), .CLK(CK), .Q(g3007), 
        .QN(n1866) );
  SDFFX1 DFF_54_Q_reg ( .D(n1885), .SI(g3007), .SE(test_se), .CLK(CK), .Q(
        test_so1), .QN() );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(test_se), .CLK(CK), .Q(
        g829), .QN(n1651) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(test_se), .CLK(CK), .Q(g1095), .QN() );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(test_se), .CLK(CK), .Q(g704), .QN() );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(test_se), .CLK(CK), .Q(g1265), .QN() );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(test_se), .CLK(CK), .Q(
        g1786), .QN() );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(test_se), .CLK(CK), .Q(g682), .QN() );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(test_se), .CLK(CK), .Q(g1296), .QN() );
  SDFFX1 DFF_62_Q_reg ( .D(g6284), .SI(g1296), .SE(test_se), .CLK(CK), .Q(
        g2602), .QN() );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(test_se), .CLK(CK), .Q(
        g8977), .QN(n1668) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(test_se), .CLK(CK), .Q(
        n3062), .QN(n1595) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(test_se), .CLK(CK), .Q(g327), 
        .QN() );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(test_se), .CLK(CK), .Q(g1389), .QN(n1603) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(test_se), .CLK(CK), .Q(
        g1371), .QN() );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(test_se), .CLK(CK), .Q(
        g1956), .QN() );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(test_se), .CLK(CK), .Q(
        g1675), .QN() );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(test_se), .CLK(CK), .Q(
        g354), .QN() );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(test_se), .CLK(CK), .Q(g113), 
        .QN() );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(test_se), .CLK(CK), .Q(g639), 
        .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(test_se), .CLK(CK), .Q(
        g1684), .QN() );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(test_se), .CLK(CK), .Q(
        g1639), .QN() );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(test_se), .CLK(CK), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(test_se), .CLK(CK), .Q(g248), .QN(n1598) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(test_se), .CLK(CK), .Q(g1707), .QN() );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(test_se), .CLK(CK), .Q(
        g1759), .QN() );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(test_se), .CLK(CK), .Q(
        g351), .QN() );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(test_se), .CLK(CK), .Q(g1957), .QN() );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(test_se), .CLK(CK), .Q(
        g1604), .QN() );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(test_se), .CLK(CK), .Q(
        g1098), .QN() );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(test_se), .CLK(CK), .Q(g932), .QN(n1591) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(test_se), .CLK(CK), .Q(g1896), .QN() );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(test_se), .CLK(CK), .Q(g736), .QN() );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(test_se), .CLK(CK), .Q(g1019), .QN() );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(test_se), .CLK(CK), .Q(
        n3061), .QN(n1625) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(test_se), .CLK(CK), .Q(g745), 
        .QN() );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(test_se), .CLK(CK), .Q(g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(test_se), .CLK(CK), .Q(
        g8979), .QN(n1667) );
  SDFFX1 DFF_92_Q_reg ( .D(n542), .SI(g8979), .SE(test_se), .CLK(CK), .Q(g32), 
        .QN() );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(test_se), .CLK(CK), .Q(n1865), 
        .QN() );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(test_se), .CLK(CK), .Q(
        g1086), .QN() );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(test_se), .CLK(CK), .Q(
        g1486), .QN() );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(test_se), .CLK(CK), .Q(
        g1730), .QN() );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(test_se), .CLK(CK), .Q(
        g1504), .QN() );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(test_se), .CLK(CK), .Q(
        g1470), .QN() );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(test_se), .CLK(CK), .Q(g822), .QN() );
  SDFFX1 DFF_100_Q_reg ( .D(g6253), .SI(g822), .SE(test_se), .CLK(CK), .Q(
        g2609), .QN() );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(test_se), .CLK(CK), .Q(
        g1678), .QN() );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(test_se), .CLK(CK), .Q(
        g174), .QN() );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(test_se), .CLK(CK), .Q(
        g1766), .QN() );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(test_se), .CLK(CK), .Q(
        g1801), .QN() );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(test_se), .CLK(CK), .Q(
        g186), .QN() );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(test_se), .CLK(CK), .Q(
        g959), .QN() );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(test_se), .CLK(CK), .Q(
        test_so2), .QN(n1869) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(test_se), .CLK(CK), .Q(
        g1407), .QN() );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(test_se), .CLK(CK), .Q(
        g1868), .QN() );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(test_se), .CLK(CK), .Q(
        g4173), .QN() );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(test_se), .CLK(CK), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(test_se), .CLK(CK), .Q(
        g396), .QN() );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(test_se), .CLK(CK), .Q(
        g1015), .QN() );
  SDFFX1 DFF_116_Q_reg ( .D(g10726), .SI(g1015), .SE(test_se), .CLK(CK), .Q(
        n1650), .QN() );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(test_se), .CLK(CK), .Q(
        n3059), .QN(n1874) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(test_se), .CLK(CK), .Q(
        g1415), .QN() );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(test_se), .CLK(CK), .Q(
        g1227), .QN() );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(test_se), .CLK(CK), .Q(
        g1721), .QN() );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(test_se), .CLK(CK), .Q(
        n3058), .QN(DFF_121_n1) );
  SDFFX1 DFF_122_Q_reg ( .D(n711), .SI(n3058), .SE(test_se), .CLK(CK), .Q(
        n3057), .QN(DFF_122_n1) );
  SDFFX1 DFF_123_Q_reg ( .D(g6934), .SI(n3057), .SE(test_se), .CLK(CK), .Q(
        g284), .QN() );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(test_se), .CLK(CK), .Q(
        g426), .QN() );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(test_se), .CLK(CK), .Q(g219), .QN() );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(test_se), .CLK(CK), .Q(
        n3056), .QN(DFF_126_n1) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(test_se), .CLK(CK), .Q(
        g806), .QN() );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(test_se), .CLK(CK), .Q(
        g1428), .QN() );
  SDFFX1 DFF_129_Q_reg ( .D(g6282), .SI(g1428), .SE(test_se), .CLK(CK), .Q(
        g2605), .QN() );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(test_se), .CLK(CK), .Q(
        g1564), .QN() );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(test_se), .CLK(CK), .Q(
        g1741), .QN(n1633) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(test_se), .CLK(CK), .Q(
        g225), .QN() );
  SDFFX1 DFF_133_Q_reg ( .D(g6928), .SI(g225), .SE(test_se), .CLK(CK), .Q(g281), .QN() );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(test_se), .CLK(CK), .Q(
        g1308), .QN() );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(test_se), .CLK(CK), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(test_se), .CLK(CK), .Q(
        n3055), .QN(DFF_136_n1) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(test_se), .CLK(CK), .Q(
        g1217), .QN() );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(test_se), .CLK(CK), .Q(
        g1589), .QN() );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(test_se), .CLK(CK), .Q(
        g1466), .QN() );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(test_se), .CLK(CK), .Q(
        g1571), .QN() );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(test_se), .CLK(CK), .Q(
        g1861), .QN() );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(test_se), .CLK(CK), .Q(
        n3054), .QN(n1688) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(test_se), .CLK(CK), .Q(
        g1448), .QN() );
  SDFFX1 DFF_145_Q_reg ( .D(g4480), .SI(g1448), .SE(test_se), .CLK(CK), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(test_se), .CLK(CK), .Q(
        g1333), .QN() );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(test_se), .CLK(CK), .Q(
        g153), .QN() );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(test_se), .CLK(CK), .Q(
        g962), .QN(n1638) );
  SDFFX1 DFF_149_Q_reg ( .D(g5536), .SI(g962), .SE(test_se), .CLK(CK), .Q(
        g4175), .QN() );
  SDFFX1 DFF_150_Q_reg ( .D(g6285), .SI(g4175), .SE(test_se), .CLK(CK), .Q(
        g2603), .QN() );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(test_se), .CLK(CK), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(test_se), .CLK(CK), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(test_se), .CLK(CK), .Q(
        g1397), .QN(n1711) );
  SDFFX1 DFF_154_Q_reg ( .D(g6283), .SI(g1397), .SE(test_se), .CLK(CK), .Q(
        g2606), .QN() );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(test_se), .CLK(CK), .Q(
        g1950), .QN() );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(test_se), .CLK(CK), .Q(g756), .QN() );
  SDFFX1 DFF_157_Q_reg ( .D(g4892), .SI(g756), .SE(test_se), .CLK(CK), .Q(
        n3053), .QN(DFF_157_n1) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(test_se), .CLK(CK), .Q(
        g549), .QN() );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(test_se), .CLK(CK), .Q(
        g105), .QN() );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(test_se), .CLK(CK), .Q(
        g1669), .QN() );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(test_se), .CLK(CK), .Q(
        test_so3), .QN() );
  SDFFX1 DFF_164_Q_reg ( .D(g6528), .SI(test_si4), .SE(test_se), .CLK(CK), .Q(
        g1531), .QN(n1652) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(test_se), .CLK(CK), .Q(
        g1458), .QN(n1703) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(test_se), .CLK(CK), .Q(
        g572), .QN() );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(test_se), .CLK(CK), .Q(
        g1011), .QN() );
  SDFFX1 DFF_168_Q_reg ( .D(g10719), .SI(g1011), .SE(test_se), .CLK(CK), .Q(
        n3051), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(test_se), .CLK(CK), .Q(
        g1411), .QN() );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(test_se), .CLK(CK), .Q(
        g1074), .QN() );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(test_se), .CLK(CK), .Q(
        g444), .QN() );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(test_se), .CLK(CK), .Q(
        g1474), .QN() );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(test_se), .CLK(CK), .Q(
        g1080), .QN() );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(test_se), .CLK(CK), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(test_se), .CLK(CK), .Q(g333), .QN() );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(test_se), .CLK(CK), .Q(g269), .QN() );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(test_se), .CLK(CK), .Q(
        g401), .QN() );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(test_se), .CLK(CK), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(test_se), .CLK(CK), .Q(g9), 
        .QN() );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(test_se), .CLK(CK), .Q(g664), 
        .QN() );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(test_se), .CLK(CK), .Q(
        g965), .QN(n1639) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(test_se), .CLK(CK), .Q(
        g1400), .QN(n1629) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(test_se), .CLK(CK), .Q(g309), .QN() );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(test_se), .CLK(CK), .Q(g814), .QN() );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(test_se), .CLK(CK), .Q(g231), .QN() );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(test_se), .CLK(CK), .Q(
        g557), .QN() );
  SDFFX1 DFF_187_Q_reg ( .D(g6283), .SI(g557), .SE(test_se), .CLK(CK), .Q(
        g2612), .QN() );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(test_se), .CLK(CK), .Q(g869), .QN() );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(test_se), .CLK(CK), .Q(
        g1383), .QN() );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(test_se), .CLK(CK), .Q(
        g158), .QN() );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(test_se), .CLK(CK), .Q(g627), .QN(n1701) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(test_se), .CLK(CK), .Q(
        g1023), .QN() );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(test_se), .CLK(CK), .Q(
        g259), .QN() );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(test_se), .CLK(CK), .Q(
        n3050), .QN(DFF_194_n1) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(test_se), .CLK(CK), .Q(
        g1327), .QN() );
  SDFFX1 DFF_196_Q_reg ( .D(g7660), .SI(g1327), .SE(test_se), .CLK(CK), .Q(
        g654), .QN() );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(test_se), .CLK(CK), .Q(g293), .QN() );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(test_se), .CLK(CK), .Q(
        g1346), .QN() );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(test_se), .CLK(CK), .Q(
        g1633), .QN() );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(test_se), .CLK(CK), .Q(
        g1753), .QN() );
  SDFFX1 DFF_201_Q_reg ( .D(n518), .SI(g1753), .SE(test_se), .CLK(CK), .Q(
        g1508), .QN(n1707) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(test_se), .CLK(CK), .Q(
        g1240), .QN() );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(test_se), .CLK(CK), .Q(
        g538), .QN() );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(test_se), .CLK(CK), .Q(
        g416), .QN() );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(test_se), .CLK(CK), .Q(
        g542), .QN() );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(test_se), .CLK(CK), .Q(
        g1681), .QN() );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(test_se), .CLK(CK), .Q(
        g374), .QN() );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(test_se), .CLK(CK), .Q(
        g563), .QN() );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(test_se), .CLK(CK), .Q(
        g1914), .QN() );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(test_se), .CLK(CK), .Q(
        g530), .QN() );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(test_se), .CLK(CK), .Q(
        g575), .QN() );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(test_se), .CLK(CK), .Q(
        g1936), .QN(n1694) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(test_se), .CLK(CK), .Q(
        g8978), .QN(n1674) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(test_se), .CLK(CK), .Q(
        test_so4), .QN(n1661) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(test_se), .CLK(CK), .Q(
        g1317), .QN() );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(test_se), .CLK(CK), .Q(
        g357), .QN() );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(test_se), .CLK(CK), .Q(
        g386), .QN() );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(test_se), .CLK(CK), .Q(
        g1601), .QN() );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(test_se), .CLK(CK), .Q(
        g166), .QN() );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(test_se), .CLK(CK), .Q(
        g501), .QN(n1690) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(test_se), .CLK(CK), .Q(g262), .QN() );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(test_se), .CLK(CK), .Q(
        g1840), .QN() );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(test_se), .CLK(CK), .Q(
        g8983), .QN(n1666) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(test_se), .CLK(CK), .Q(g318), .QN() );
  SDFFX1 DFF_226_Q_reg ( .D(g5763), .SI(g318), .SE(test_se), .CLK(CK), .Q(
        g1356), .QN() );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(test_se), .CLK(CK), .Q(
        g794), .QN() );
  SDFFX1 DFF_228_Q_reg ( .D(g10722), .SI(g794), .SE(test_se), .CLK(CK), .Q(
        n3048), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(test_se), .CLK(CK), .Q(
        g302), .QN() );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(test_se), .CLK(CK), .Q(
        g342), .QN() );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(test_se), .CLK(CK), .Q(
        g1250), .QN() );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(test_se), .CLK(CK), .Q(
        g1163), .QN() );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(test_se), .CLK(CK), .Q(
        n3047), .QN(g8271) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(test_se), .CLK(CK), .Q(
        g1032), .QN() );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(test_se), .CLK(CK), .Q(
        g1432), .QN() );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(test_se), .CLK(CK), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(test_se), .CLK(CK), .Q(
        g363), .QN() );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(test_se), .CLK(CK), .Q(g330), 
        .QN() );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(test_se), .CLK(CK), .Q(
        g1157), .QN() );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(test_se), .CLK(CK), .Q(
        n3046), .QN(n1648) );
  SDFFX1 DFF_242_Q_reg ( .D(g10721), .SI(n3046), .SE(test_se), .CLK(CK), .Q(
        n3045), .QN(DFF_242_n1) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(test_se), .CLK(CK), .Q(
        g928), .QN(n1604) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(test_se), .CLK(CK), .Q(g261), .QN() );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(test_se), .CLK(CK), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(test_se), .CLK(CK), .Q(g254), .QN() );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(test_se), .CLK(CK), .Q(
        g4178), .QN() );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(test_se), .CLK(CK), .Q(g861), .QN() );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(test_se), .CLK(CK), .Q(
        g1627), .QN() );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(test_se), .CLK(CK), .Q(
        g1292), .QN() );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(test_se), .CLK(CK), .Q(
        g290), .QN() );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(test_se), .CLK(CK), .Q(
        n3044), .QN(n1873) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(test_se), .CLK(CK), .Q(
        g4176), .QN() );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(test_se), .CLK(CK), .Q(
        g1583), .QN() );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(test_se), .CLK(CK), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(test_se), .CLK(CK), .Q(
        g1561), .QN() );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(test_se), .CLK(CK), .Q(
        g1546), .QN() );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(test_se), .CLK(CK), .Q(
        g287), .QN() );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(test_se), .CLK(CK), .Q(
        g560), .QN() );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(test_se), .CLK(CK), .Q(g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n667), .SI(g617), .SE(test_se), .CLK(CK), .Q(n1631), .QN() );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(test_se), .CLK(CK), .Q(
        g336), .QN() );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(test_se), .CLK(CK), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(test_se), .CLK(CK), .Q(g305), 
        .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(test_se), .CLK(CK), .Q(
        g345), .QN() );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(test_se), .CLK(CK), .Q(g8), 
        .QN() );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(test_se), .CLK(CK), .Q(
        test_so5), .QN() );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(test_se), .CLK(CK), .Q(
        g2648), .QN() );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(test_se), .CLK(CK), .Q(
        g255), .QN() );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(test_se), .CLK(CK), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(test_se), .CLK(CK), .Q(
        g1738), .QN(n1640) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(test_se), .CLK(CK), .Q(
        g1478), .QN() );
  SDFFX1 DFF_275_Q_reg ( .D(n562), .SI(g1478), .SE(test_se), .CLK(CK), .Q(
        n3042), .QN(DFF_275_n1) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(test_se), .CLK(CK), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(test_se), .CLK(CK), .Q(
        g1482), .QN() );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(test_se), .CLK(CK), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(test_se), .CLK(CK), .Q(
        g296), .QN() );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(test_se), .CLK(CK), .Q(
        g1663), .QN() );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(test_se), .CLK(CK), .Q(
        g700), .QN() );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(test_se), .CLK(CK), .Q(
        g1762), .QN() );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(test_se), .CLK(CK), .Q(
        g360), .QN() );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(test_se), .CLK(CK), .Q(g192), .QN() );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(test_se), .CLK(CK), .Q(
        g1657), .QN() );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(test_se), .CLK(CK), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(test_se), .CLK(CK), .Q(
        g8980), .QN(n1673) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(test_se), .CLK(CK), .Q(
        g566), .QN() );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(test_se), .CLK(CK), .Q(
        n3041), .QN(n1714) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(test_se), .CLK(CK), .Q(
        g1089), .QN() );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(test_se), .CLK(CK), .Q(
        g2986), .QN() );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(test_se), .CLK(CK), .Q(
        g1071), .QN() );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(test_se), .CLK(CK), .Q(
        g986), .QN(n1722) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(test_se), .CLK(CK), .Q(
        g971), .QN() );
  SDFFX1 DFF_295_Q_reg ( .D(g6265), .SI(g971), .SE(test_se), .CLK(CK), .Q(
        g1955), .QN() );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(test_se), .CLK(CK), .Q(
        g143), .QN() );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(test_se), .CLK(CK), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(test_se), .CLK(CK), .Q(
        g1212), .QN() );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(test_se), .CLK(CK), .Q(
        g1918), .QN() );
  SDFFX1 DFF_301_Q_reg ( .D(g7705), .SI(g1918), .SE(test_se), .CLK(CK), .Q(
        g4179), .QN() );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(test_se), .CLK(CK), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(test_se), .CLK(CK), .Q(
        g237), .QN() );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(test_se), .CLK(CK), .Q(g746), 
        .QN() );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(test_se), .CLK(CK), .Q(
        g1462), .QN() );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(test_se), .CLK(CK), .Q(
        g178), .QN() );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(test_se), .CLK(CK), .Q(
        g366), .QN() );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(test_se), .CLK(CK), .Q(g837), 
        .QN() );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(test_se), .CLK(CK), .Q(g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(test_se), .CLK(CK), .Q(
        g1854), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(test_se), .CLK(CK), .Q(
        g944), .QN() );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(test_se), .CLK(CK), .Q(
        g1941), .QN() );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(test_se), .CLK(CK), .Q(
        g170), .QN() );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(test_se), .CLK(CK), .Q(
        g1520), .QN(n1710) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(test_se), .CLK(CK), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(test_se), .CLK(CK), .Q(
        g953), .QN() );
  SDFFX1 DFF_318_Q_reg ( .D(g5556), .SI(g953), .SE(test_se), .CLK(CK), .Q(
        g1958), .QN() );
  SDFFX1 DFF_319_Q_reg ( .D(g10664), .SI(g1958), .SE(test_se), .CLK(CK), .Q(
        n3040), .QN(DFF_319_n1) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(test_se), .CLK(CK), .Q(
        g1765), .QN() );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(test_se), .CLK(CK), .Q(
        g1733), .QN() );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(test_se), .CLK(CK), .Q(
        test_so6), .QN() );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(test_se), .CLK(CK), .Q(
        g1610), .QN() );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(test_se), .CLK(CK), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(test_se), .CLK(CK), .Q(
        g1324), .QN() );
  SDFFX1 DFF_326_Q_reg ( .D(g6541), .SI(g1324), .SE(test_se), .CLK(CK), .Q(
        g1540), .QN() );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(test_se), .CLK(CK), .Q(
        n3038), .QN(n1624) );
  SDFFX1 DFF_328_Q_reg ( .D(n687), .SI(n3038), .SE(test_se), .CLK(CK), .Q(
        g3069), .QN() );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(test_se), .CLK(CK), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(test_se), .CLK(CK), .Q(
        n3037), .QN(DFF_330_n1) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(test_se), .CLK(CK), .Q(
        g213), .QN() );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(test_se), .CLK(CK), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(test_se), .CLK(CK), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(test_se), .CLK(CK), .Q(
        g1245), .QN() );
  SDFFX1 DFF_335_Q_reg ( .D(n550), .SI(g1245), .SE(test_se), .CLK(CK), .Q(
        n3036), .QN(n1683) );
  SDFFX1 DFF_336_Q_reg ( .D(g6672), .SI(n3036), .SE(test_se), .CLK(CK), .Q(
        n3035), .QN(DFF_336_n1) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(test_se), .CLK(CK), .Q(
        g148), .QN() );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(test_se), .CLK(CK), .Q(g833), 
        .QN() );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(test_se), .CLK(CK), .Q(
        g1923), .QN(n1718) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(test_se), .CLK(CK), .Q(
        g936), .QN(n1630) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(test_se), .CLK(CK), .Q(
        g1314), .QN() );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(test_se), .CLK(CK), .Q(g849), .QN() );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(test_se), .CLK(CK), .Q(
        g1336), .QN() );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(test_se), .CLK(CK), .Q(
        g272), .QN() );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(test_se), .CLK(CK), .Q(
        g1806), .QN() );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(test_se), .CLK(CK), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(test_se), .CLK(CK), .Q(
        g1887), .QN() );
  SDFFX1 DFF_350_Q_reg ( .D(g10724), .SI(g1887), .SE(test_se), .CLK(CK), .Q(
        n3034), .QN(DFF_350_n1) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(test_se), .CLK(CK), .Q(
        g968), .QN() );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(test_se), .CLK(CK), .Q(
        n3033), .QN(n1642) );
  SDFFX1 DFF_353_Q_reg ( .D(g4484), .SI(n3033), .SE(test_se), .CLK(CK), .Q(
        g1137), .QN(n1597) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(test_se), .CLK(CK), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(test_se), .CLK(CK), .Q(
        g1255), .QN() );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(test_se), .CLK(CK), .Q(
        g257), .QN() );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(test_se), .CLK(CK), .Q(g874), .QN() );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(test_se), .CLK(CK), .Q(g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(test_se), .CLK(CK), .Q(g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(test_se), .CLK(CK), .Q(g636), .QN() );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(test_se), .CLK(CK), .Q(
        g1218), .QN() );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(test_se), .CLK(CK), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(test_se), .CLK(CK), .Q(
        g8986), .QN(n1665) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(test_se), .CLK(CK), .Q(
        g182), .QN() );
  SDFFX1 DFF_365_Q_reg ( .D(g11303), .SI(g182), .SE(test_se), .CLK(CK), .Q(
        g950), .QN() );
  SDFFX1 DFF_366_Q_reg ( .D(g4477), .SI(g950), .SE(test_se), .CLK(CK), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(test_se), .CLK(CK), .Q(g857), .QN() );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(test_se), .CLK(CK), .Q(
        g448), .QN() );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(test_se), .CLK(CK), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(test_se), .CLK(CK), .Q(
        g1727), .QN() );
  SDFFX1 DFF_371_Q_reg ( .D(g6470), .SI(g1727), .SE(test_se), .CLK(CK), .Q(
        g1592), .QN() );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(test_se), .CLK(CK), .Q(
        g1703), .QN() );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(test_se), .CLK(CK), .Q(
        g1932), .QN() );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(test_se), .CLK(CK), .Q(
        g1624), .QN() );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(test_se), .CLK(CK), .Q(
        test_so7), .QN() );
  SDFFX1 DFF_377_Q_reg ( .D(g6281), .SI(test_si8), .SE(test_se), .CLK(CK), .Q(
        g2601), .QN() );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(test_se), .CLK(CK), .Q(
        g440), .QN() );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(test_se), .CLK(CK), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(test_se), .CLK(CK), .Q(g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(test_se), .CLK(CK), .Q(g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(test_se), .CLK(CK), .Q(g139), .QN() );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(test_se), .CLK(CK), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(g10720), .SI(g1149), .SE(test_se), .CLK(CK), .Q(
        n3031), .QN(DFF_384_n1) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(test_se), .CLK(CK), .Q(
        n3030), .QN(DFF_385_n1) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(test_se), .CLK(CK), .Q(
        g263), .QN() );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(test_se), .CLK(CK), .Q(g818), .QN() );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(test_se), .CLK(CK), .Q(
        g1747), .QN() );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(test_se), .CLK(CK), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(test_se), .CLK(CK), .Q(g275), .QN() );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(test_se), .CLK(CK), .Q(
        g1524), .QN(n1649) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(test_se), .CLK(CK), .Q(
        g1577), .QN() );
  SDFFX1 DFF_393_Q_reg ( .D(g6733), .SI(g1577), .SE(test_se), .CLK(CK), .Q(
        g810), .QN() );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(test_se), .CLK(CK), .Q(
        g391), .QN() );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(test_se), .CLK(CK), .Q(g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(test_se), .CLK(CK), .Q(
        g1386), .QN() );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(test_se), .CLK(CK), .Q(
        g253), .QN() );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(test_se), .CLK(CK), .Q(g875), .QN() );
  SDFFX1 DFF_399_Q_reg ( .D(g4473), .SI(g875), .SE(test_se), .CLK(CK), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(test_se), .CLK(CK), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(test_se), .CLK(CK), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(test_se), .CLK(CK), .Q(
        g1083), .QN() );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(test_se), .CLK(CK), .Q(
        g650), .QN(n1709) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(test_se), .CLK(CK), .Q(
        g1636), .QN() );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(test_se), .CLK(CK), .Q(g853), .QN() );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(test_se), .CLK(CK), .Q(
        g421), .QN() );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(test_se), .CLK(CK), .Q(
        g4174), .QN() );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(test_se), .CLK(CK), .Q(
        g956), .QN() );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(test_se), .CLK(CK), .Q(
        g378), .QN() );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(test_se), .CLK(CK), .Q(
        g1756), .QN() );
  SDFFX1 DFF_411_Q_reg ( .D(g6253), .SI(g1756), .SE(test_se), .CLK(CK), .Q(
        g2604), .QN() );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(test_se), .CLK(CK), .Q(g841), .QN() );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(test_se), .CLK(CK), .Q(
        g1027), .QN() );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(test_se), .CLK(CK), .Q(
        g1003), .QN() );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(test_se), .CLK(CK), .Q(
        g1403), .QN() );
  SDFFX1 DFF_416_Q_reg ( .D(g4498), .SI(g1403), .SE(test_se), .CLK(CK), .Q(
        g1145), .QN(n1617) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(test_se), .CLK(CK), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(test_se), .CLK(CK), .Q(
        g1223), .QN() );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(test_se), .CLK(CK), .Q(
        g406), .QN() );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(test_se), .CLK(CK), .Q(
        g1811), .QN(n1699) );
  SDFFX1 DFF_421_Q_reg ( .D(g10784), .SI(g1811), .SE(test_se), .CLK(CK), .Q(
        n3029), .QN(n1684) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(test_se), .CLK(CK), .Q(
        g1654), .QN() );
  SDFFX1 DFF_424_Q_reg ( .D(g6332), .SI(g1654), .SE(test_se), .CLK(CK), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(test_se), .CLK(CK), .Q(
        g1595), .QN() );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(test_se), .CLK(CK), .Q(
        g1537), .QN(n1636) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(test_se), .CLK(CK), .Q(
        g727), .QN() );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(test_se), .CLK(CK), .Q(
        test_so8), .QN() );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(test_se), .CLK(CK), .Q(
        g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(test_se), .CLK(CK), .Q(
        g481), .QN(n1680) );
  SDFFX1 DFF_431_Q_reg ( .D(g3462), .SI(g481), .SE(test_se), .CLK(CK), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(test_se), .CLK(CK), .Q(
        g1330), .QN() );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(test_se), .CLK(CK), .Q(g845), .QN() );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(test_se), .CLK(CK), .Q(
        g4181), .QN() );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(test_se), .CLK(CK), .Q(
        g1512), .QN() );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(test_se), .CLK(CK), .Q(
        n3027), .QN(DFF_436_n1) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(test_se), .CLK(CK), .Q(
        g1490), .QN() );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(test_se), .CLK(CK), .Q(
        g1166), .QN() );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(test_se), .CLK(CK), .Q(
        g348), .QN() );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(test_se), .CLK(CK), .Q(n3026), .QN(DFF_441_n1) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(test_se), .CLK(CK), .Q(
        g1260), .QN() );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(test_se), .CLK(CK), .Q(
        g260), .QN() );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(test_se), .CLK(CK), .Q(g131), .QN() );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(test_se), .CLK(CK), .Q(
        n3025), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(test_se), .CLK(CK), .Q(
        g258), .QN() );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(test_se), .CLK(CK), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(test_se), .CLK(CK), .Q(
        g1318), .QN() );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(test_se), .CLK(CK), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(test_se), .CLK(CK), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g6285), .SI(g677), .SE(test_se), .CLK(CK), .Q(
        g2608), .QN() );
  SDFFX1 DFF_452_Q_reg ( .D(n519), .SI(g2608), .SE(test_se), .CLK(CK), .Q(
        n3024), .QN(DFF_452_n1) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(test_se), .CLK(CK), .Q(
        g1549), .QN() );
  SDFFX1 DFF_454_Q_reg ( .D(g11300), .SI(g1549), .SE(test_se), .CLK(CK), .Q(
        g947), .QN() );
  SDFFX1 DFF_455_Q_reg ( .D(g9555), .SI(g947), .SE(test_se), .CLK(CK), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(test_se), .CLK(CK), .Q(
        g1598), .QN() );
  SDFFX1 DFF_457_Q_reg ( .D(g4471), .SI(g1598), .SE(test_se), .CLK(CK), .Q(
        g1121), .QN(n1618) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(test_se), .CLK(CK), .Q(
        g1321), .QN() );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(test_se), .CLK(CK), .Q(
        g506), .QN(n1600) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(test_se), .CLK(CK), .Q(
        g546), .QN() );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(test_se), .CLK(CK), .Q(
        g1909), .QN() );
  SDFFX1 DFF_462_Q_reg ( .D(g6265), .SI(g1909), .SE(test_se), .CLK(CK), .Q(
        g755), .QN() );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(test_se), .CLK(CK), .Q(
        g1552), .QN() );
  SDFFX1 DFF_464_Q_reg ( .D(g6281), .SI(g1552), .SE(test_se), .CLK(CK), .Q(
        g2610), .QN() );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(test_se), .CLK(CK), .Q(
        g1687), .QN() );
  SDFFX1 DFF_466_Q_reg ( .D(g6514), .SI(g1687), .SE(test_se), .CLK(CK), .Q(
        g1586), .QN() );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(test_se), .CLK(CK), .Q(g324), .QN() );
  SDFFX1 DFF_468_Q_reg ( .D(g4490), .SI(g324), .SE(test_se), .CLK(CK), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(test_se), .CLK(CK), .Q(
        g1341), .QN() );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(test_se), .CLK(CK), .Q(
        g1710), .QN() );
  SDFFX1 DFF_472_Q_reg ( .D(g10785), .SI(g1710), .SE(test_se), .CLK(CK), .Q(
        n3023), .QN(n1623) );
  SDFFX1 DFF_473_Q_reg ( .D(g6179), .SI(n3023), .SE(test_se), .CLK(CK), .Q(
        n3022), .QN(n1634) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(test_se), .CLK(CK), .Q(
        g135), .QN() );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(test_se), .CLK(CK), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g6284), .SI(g525), .SE(test_se), .CLK(CK), .Q(
        g2607), .QN() );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(test_se), .CLK(CK), .Q(
        g1607), .QN() );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(test_se), .CLK(CK), .Q(g321), .QN() );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(test_se), .CLK(CK), .Q(
        g8982), .QN(n1672) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(test_se), .CLK(CK), .Q(
        g1275), .QN() );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(test_se), .CLK(CK), .Q(
        test_so9), .QN() );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(test_se), .CLK(CK), 
        .Q(g1615), .QN() );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(test_se), .CLK(CK), .Q(
        g382), .QN() );
  SDFFX1 DFF_484_Q_reg ( .D(g6331), .SI(g382), .SE(test_se), .CLK(CK), .Q(
        n3020), .QN(n1700) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(test_se), .CLK(CK), .Q(
        g266), .QN() );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(test_se), .CLK(CK), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(test_se), .CLK(CK), .Q(
        n3019), .QN(n1687) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(test_se), .CLK(CK), .Q(
        g673), .QN() );
  SDFFX1 DFF_489_Q_reg ( .D(g4904), .SI(g673), .SE(test_se), .CLK(CK), .Q(
        n3018), .QN(DFF_489_n1) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(test_se), .CLK(CK), .Q(
        g162), .QN() );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(test_se), .CLK(CK), .Q(
        g411), .QN() );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(test_se), .CLK(CK), .Q(
        g431), .QN(n1876) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(test_se), .CLK(CK), .Q(
        g1905), .QN() );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(test_se), .CLK(CK), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(test_se), .CLK(CK), .Q(
        g1630), .QN() );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(test_se), .CLK(CK), .Q(
        g8976), .QN(n1671) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(test_se), .CLK(CK), .Q(
        g991), .QN(n1871) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(test_se), .CLK(CK), .Q(
        g1300), .QN() );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(test_se), .CLK(CK), .Q(
        g339), .QN() );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(test_se), .CLK(CK), .Q(g256), .QN() );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(test_se), .CLK(CK), .Q(
        g1750), .QN() );
  SDFFX1 DFF_502_Q_reg ( .D(g6282), .SI(g1750), .SE(test_se), .CLK(CK), .Q(
        g2611), .QN() );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(test_se), .CLK(CK), .Q(
        g1440), .QN() );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(test_se), .CLK(CK), .Q(
        g1666), .QN() );
  SDFFX1 DFF_505_Q_reg ( .D(g6522), .SI(g1666), .SE(test_se), .CLK(CK), .Q(
        g1528), .QN(n1635) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(test_se), .CLK(CK), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(g10780), .SI(g1351), .SE(test_se), .CLK(CK), .Q(
        n3017), .QN(n1601) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(test_se), .CLK(CK), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(test_se), .CLK(CK), .Q(
        g1618), .QN() );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(test_se), .CLK(CK), .Q(
        g1235), .QN() );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(test_se), .CLK(CK), .Q(
        g299), .QN() );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(test_se), .CLK(CK), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(test_se), .CLK(CK), .Q(
        g8981), .QN(n1664) );
  SDFFX1 DFF_514_Q_reg ( .D(g6534), .SI(g8981), .SE(test_se), .CLK(CK), .Q(
        g1555), .QN() );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(test_se), .CLK(CK), .Q(
        g995), .QN() );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(test_se), .CLK(CK), .Q(
        g1621), .QN() );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(test_se), .CLK(CK), .Q(
        n3016), .QN(n1596) );
  SDFFX1 DFF_518_Q_reg ( .D(g7441), .SI(n3016), .SE(test_se), .CLK(CK), .Q(
        g643), .QN(n1612) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(test_se), .CLK(CK), .Q(
        g1494), .QN() );
  SDFFX1 DFF_520_Q_reg ( .D(g6468), .SI(g1494), .SE(test_se), .CLK(CK), .Q(
        g1567), .QN() );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(test_se), .CLK(CK), .Q(
        g691), .QN() );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(test_se), .CLK(CK), .Q(
        g534), .QN() );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(test_se), .CLK(CK), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(test_se), .CLK(CK), .Q(
        g569), .QN() );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(test_se), .CLK(CK), .Q(
        g1160), .QN() );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(test_se), .CLK(CK), .Q(
        g1360), .QN() );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(test_se), .CLK(CK), .Q(g1), 
        .QN() );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(test_se), .CLK(CK), .Q(g511), 
        .QN(n1679) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(test_se), .CLK(CK), .Q(
        g1724), .QN() );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(test_se), .CLK(CK), .Q(g12), .QN() );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(test_se), .CLK(CK), .Q(g1878), .QN() );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(test_se), .CLK(CK), .Q(
        g8984), .QN(n1670) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(test_se), .CLK(CK), .Q(
        g1101), .QN(n1654) );
  NAND2X1 U1553 ( .A(n1173), .B(1'b1), .Q(n1169) );
  NAND2X1 U1554 ( .A(n1173), .B(1'b1), .Q(n1167) );
  NAND3X1 U1555 ( .A(n1145), .B(1'b1), .C(n1976), .Q(n1142) );
  AO222X1 U1556 ( .A(g1351), .B(n1511), .C(g4208), .D(n1512), .E(
        g1324), .F(n576), .Q(n1510) );
  AND4X1 U1557 ( .A(n1574), .B(n1578), .C(g6257), .D(g6258), .Q(n1507)
         );
  AND4X1 U1558 ( .A(n1574), .B(n1396), .C(g6260), .D(g6259), .Q(n1508)
         );
  AND2X1 U1559 ( .A(n798), .B(n1569), .Q(n1574) );
  NAND4X1 U1560 ( .A(n1569), .B(n842), .C(g6262), .D(n1570), .Q(n1541) );
  AOI222X1 U1561 ( .A(g1546), .B(n1486), .C(g4203), .D(n1481), .E(
        g1589), .F(n1485), .Q(n1555) );
  INVX1 U1562 ( .IN(n1360), .Q(n526) );
  INVX1 U1563 ( .IN(n1484), .Q(n583) );
  INVX1 U1564 ( .IN(n1899), .Q(n1891) );
  AO222X1 U1565 ( .A(g4206), .B(n1512), .C(g4197), .D(n1481), .E(
        g1341), .F(n1511), .Q(n1531) );
  AND4X1 U1566 ( .A(g6260), .B(g6259), .C(g6258), .D(n1544), .Q(n1581)
         );
  AO222X1 U1567 ( .A(g1346), .B(n1511), .C(g4207_Payload), .D(n1512), .E(
        g1321), .F(n576), .Q(n1521) );
  INVX1 U1568 ( .IN(n1889), .Q(n1904) );
  INVX1 U1569 ( .IN(n1890), .Q(n1906) );
  INVX1 U1570 ( .IN(n1898), .Q(n1892) );
  AND2X1 U1571 ( .A(n796), .B(n1569), .Q(n1544) );
  NAND3X1 U1572 ( .A(g6258), .B(n1849), .C(n1580), .Q(n1545) );
  AND2X1 U1573 ( .A(n1395), .B(n1569), .Q(n1548) );
  AO22X1 U1574 ( .A(n583), .B(n1569), .C(n1583), .D(n1833), .Q(n842)
         );
  AO22X1 U1575 ( .A(n1114), .B(n1285), .C(n1326), .D(n629), .Q(n1284)
         );
  AO221X1 U1576 ( .A(g1318), .B(n576), .C(g4209), .D(n1476), .E(
        n1531), .Q(n1527) );
  AO221X1 U1577 ( .A(g4196), .B(n1530), .C(g4192), .D(n1507), .E(
        n1509), .Q(n1528) );
  AOI22X1 U1578 ( .A(g1327), .B(n576), .C(g4212), .D(n1476), .Q(n1493) );
  AO221X1 U1579 ( .A(g4210), .B(n1476), .C(g1), .D(n578), .E(n1521), 
        .Q(n1518) );
  AO221X1 U1580 ( .A(g4193), .B(n1507), .C(g936), .D(n1508), .E(
        n1509), .Q(n1519) );
  AO221X1 U1581 ( .A(g4211), .B(n1476), .C(g8), .D(n578), .E(n1510), 
        .Q(n1503) );
  AO221X1 U1582 ( .A(g4194), .B(n1507), .C(g940), .D(n1508), .E(
        n1509), .Q(n1504) );
  AO222X1 U1583 ( .A(g4216), .B(n1512), .C(g4195), .D(n1481), .E(
        g1336), .F(n1511), .Q(n1540) );
  OA22X1 U1584 ( .A(n1420), .B(n1681), .C(n1434), .D(n625), .Q(n1390)
         );
  AOI22X1 U1585 ( .A(g1330), .B(n576), .C(g4213), .D(n1476), .Q(n1475) );
  ISOLANDX1 U1586 ( .D(n524), .ISO(n1856), .Q(n1855) );
  INVX1 U1587 ( .IN(n1855), .Q(n1361) );
  INVX1 U1588 ( .IN(n1349), .Q(n527) );
  INVX1 U1589 ( .IN(n1908), .Q(n1903) );
  NOR2X1 U1590 ( .A(n794), .B(n1464), .Q(g11206) );
  NAND2X1 U1591 ( .A(n1887), .B(n793), .Q(g10801) );
  AOI22X1 U1592 ( .A(test_so9), .B(n1511), .C(g4215), .D(n1476), .Q(
        n1551) );
  NAND2X1 U1593 ( .A(n526), .B(g369), .Q(n1389) );
  AOI222X1 U1594 ( .A(g1721), .B(n575), .C(g1314), .D(n576), .E(
        g4205), .F(n1476), .Q(n1534) );
  AOI222X1 U1595 ( .A(g4201), .B(n1481), .C(g302), .D(n1482), .E(
        g278), .F(n1483), .Q(n1469) );
  INVX1 U1596 ( .IN(n1337), .Q(n524) );
  NAND4X1 U1597 ( .A(n1440), .B(n1651), .C(n1441), .D(n1442), .Q(
        n1239) );
  NAND2X1 U1598 ( .A(g750), .B(n1647), .Q(n1592) );
  INVX1 U1599 ( .IN(g1696), .Q(n1723) );
  INVX1 U1600 ( .IN(n1723), .Q(n1724) );
  INVX1 U1601 ( .IN(g99), .Q(n1725) );
  INVX1 U1602 ( .IN(n1725), .Q(g6279) );
  INVX1 U1603 ( .IN(g96), .Q(n1727) );
  INVX1 U1604 ( .IN(n1727), .Q(g6278) );
  INVX1 U1605 ( .IN(g95), .Q(n1729) );
  INVX1 U1606 ( .IN(n1729), .Q(g6277) );
  INVX1 U1607 ( .IN(g94), .Q(n1731) );
  INVX1 U1608 ( .IN(n1731), .Q(g6276) );
  INVX1 U1609 ( .IN(g93), .Q(n1733) );
  INVX1 U1610 ( .IN(n1733), .Q(g6275) );
  INVX1 U1611 ( .IN(g92), .Q(n1735) );
  INVX1 U1612 ( .IN(n1735), .Q(g6274) );
  INVX1 U1613 ( .IN(g91), .Q(n1737) );
  INVX1 U1614 ( .IN(n1737), .Q(g6273) );
  INVX1 U1615 ( .IN(g90), .Q(n1739) );
  INVX1 U1616 ( .IN(n1739), .Q(g6272) );
  INVX1 U1617 ( .IN(g89), .Q(n1741) );
  INVX1 U1618 ( .IN(n1741), .Q(g6271) );
  INVX1 U1619 ( .IN(g88), .Q(n1743) );
  INVX1 U1620 ( .IN(n1743), .Q(g6270) );
  INVX1 U1621 ( .IN(g87), .Q(n1745) );
  INVX1 U1622 ( .IN(n1745), .Q(g6269) );
  INVX1 U1623 ( .IN(g86), .Q(n1747) );
  INVX1 U1624 ( .IN(n1747), .Q(g6268) );
  INVX1 U1625 ( .IN(g85), .Q(n1749) );
  INVX1 U1626 ( .IN(n1749), .Q(g6267) );
  INVX1 U1627 ( .IN(g84), .Q(n1751) );
  INVX1 U1628 ( .IN(n1751), .Q(g6266) );
  INVX1 U1629 ( .IN(g27), .Q(n1753) );
  INVX1 U1630 ( .IN(n1753), .Q(g7744) );
  INVX1 U1631 ( .IN(g1961), .Q(n1755) );
  INVX1 U1632 ( .IN(n1755), .Q(g4887) );
  INVX1 U1633 ( .IN(g1960), .Q(n1757) );
  INVX1 U1634 ( .IN(n1757), .Q(g4888) );
  INVX1 U1635 ( .IN(g100), .Q(n1759) );
  INVX1 U1636 ( .IN(n1759), .Q(g6280) );
  INVX1 U1637 ( .IN(g1191), .Q(n1761) );
  INVX1 U1638 ( .IN(n1761), .Q(g4215) );
  INVX1 U1639 ( .IN(g1185), .Q(n1763) );
  INVX1 U1640 ( .IN(n1763), .Q(g4213) );
  INVX1 U1641 ( .IN(g1182), .Q(n1765) );
  INVX1 U1642 ( .IN(n1765), .Q(g4212) );
  INVX1 U1643 ( .IN(g910), .Q(n1767) );
  INVX1 U1644 ( .IN(n1767), .Q(g4200) );
  INVX1 U1645 ( .IN(g916), .Q(n1769) );
  INVX1 U1646 ( .IN(n1769), .Q(g4202) );
  INVX1 U1647 ( .IN(g913), .Q(n1771) );
  INVX1 U1648 ( .IN(n1771), .Q(g4201) );
  INVX1 U1649 ( .IN(g82), .Q(n1773) );
  INVX1 U1650 ( .IN(n1773), .Q(g6264) );
  INVX1 U1651 ( .IN(g31), .Q(n1775) );
  INVX1 U1652 ( .IN(n1775), .Q(g6255) );
  INVX1 U1653 ( .IN(g1170), .Q(n1777) );
  INVX1 U1654 ( .IN(n1777), .Q(g4205) );
  INVX1 U1655 ( .IN(g919), .Q(n1779) );
  INVX1 U1656 ( .IN(n1779), .Q(g4203) );
  INVX1 U1657 ( .IN(g907), .Q(n1781) );
  INVX1 U1658 ( .IN(n1781), .Q(g4199) );
  INVX1 U1659 ( .IN(g904), .Q(n1783) );
  INVX1 U1660 ( .IN(n1783), .Q(g4198) );
  INVX1 U1661 ( .IN(g886), .Q(n1785) );
  INVX1 U1662 ( .IN(n1785), .Q(g4191) );
  INVX1 U1663 ( .IN(g1188), .Q(n1787) );
  INVX1 U1664 ( .IN(n1787), .Q(g4214) );
  INVX1 U1665 ( .IN(g889), .Q(n1789) );
  INVX1 U1666 ( .IN(n1789), .Q(g4192) );
  INVX1 U1667 ( .IN(g1173), .Q(n1791) );
  INVX1 U1668 ( .IN(n1791), .Q(g4209) );
  INVX1 U1669 ( .IN(g922), .Q(n1793) );
  INVX1 U1670 ( .IN(n1793), .Q(g4204) );
  INVX1 U1671 ( .IN(g901), .Q(n1795) );
  INVX1 U1672 ( .IN(n1795), .Q(g4197) );
  INVX1 U1673 ( .IN(g898), .Q(n1797) );
  INVX1 U1674 ( .IN(n1797), .Q(g4195) );
  INVX1 U1675 ( .IN(g1203), .Q(n1799) );
  INVX1 U1676 ( .IN(n1799), .Q(g4208) );
  INVX1 U1677 ( .IN(g1200), .Q(n1801) );
  INVX1 U1678 ( .IN(n1801), .Q(g4207_Payload) );
  INVX1 U1679 ( .IN(g1197), .Q(n1803) );
  INVX1 U1680 ( .IN(n1803), .Q(g4206) );
  INVX1 U1681 ( .IN(g1194), .Q(n1805) );
  INVX1 U1682 ( .IN(n1805), .Q(g4216) );
  INVX1 U1683 ( .IN(g925), .Q(n1807) );
  INVX1 U1684 ( .IN(n1807), .Q(g4196) );
  INVX1 U1685 ( .IN(g895), .Q(n1809) );
  INVX1 U1686 ( .IN(n1809), .Q(g4194) );
  INVX1 U1687 ( .IN(g892), .Q(n1811) );
  INVX1 U1688 ( .IN(n1811), .Q(g4193) );
  INVX1 U1689 ( .IN(g1179), .Q(n1813) );
  INVX1 U1690 ( .IN(n1813), .Q(g4211) );
  INVX1 U1691 ( .IN(g1176), .Q(n1815) );
  INVX1 U1692 ( .IN(n1815), .Q(g4210) );
  INVX1 U1693 ( .IN(g83), .Q(n1817) );
  INVX1 U1694 ( .IN(n1817), .Q(g6265) );
  INVX1 U1695 ( .IN(g29), .Q(n1819) );
  INVX1 U1696 ( .IN(n1819), .Q(g6253) );
  INVX1 U1697 ( .IN(g28), .Q(n1821) );
  INVX1 U1698 ( .IN(n1821), .Q(g6285) );
  INVX1 U1699 ( .IN(g104), .Q(n1823) );
  INVX1 U1700 ( .IN(n1823), .Q(g6284) );
  INVX1 U1701 ( .IN(g103), .Q(n1825) );
  INVX1 U1702 ( .IN(n1825), .Q(g6283) );
  INVX1 U1703 ( .IN(g102), .Q(n1827) );
  INVX1 U1704 ( .IN(n1827), .Q(g6282) );
  INVX1 U1705 ( .IN(g101), .Q(n1829) );
  INVX1 U1706 ( .IN(n1829), .Q(g6281) );
  INVX1 U1707 ( .IN(g46), .Q(n1831) );
  INVX1 U1708 ( .IN(n1831), .Q(g6261) );
  INVX1 U1709 ( .IN(g30), .Q(n1833) );
  INVX1 U1710 ( .IN(n1833), .Q(g6254) );
  INVX1 U1711 ( .IN(g41), .Q(n1835) );
  INVX1 U1712 ( .IN(n1835), .Q(g6256) );
  INVX1 U1713 ( .IN(g873), .Q(n1837) );
  INVX1 U1714 ( .IN(n1837), .Q(g5105) );
  INVX1 U1715 ( .IN(g872), .Q(n1839) );
  INVX1 U1716 ( .IN(n1839), .Q(g5101) );
  INVX1 U1717 ( .IN(g47), .Q(n1841) );
  INVX1 U1718 ( .IN(n1841), .Q(g6262) );
  INVX1 U1719 ( .IN(g48), .Q(n1843) );
  INVX1 U1720 ( .IN(n1843), .Q(g6263) );
  INVX1 U1721 ( .IN(g45), .Q(n1845) );
  INVX1 U1722 ( .IN(n1845), .Q(g6260) );
  INVX1 U1723 ( .IN(g44), .Q(n1847) );
  INVX1 U1724 ( .IN(n1847), .Q(g6259) );
  INVX1 U1725 ( .IN(g42), .Q(n1849) );
  INVX1 U1726 ( .IN(n1849), .Q(g6257) );
  INVX1 U1727 ( .IN(g43), .Q(n1851) );
  INVX1 U1728 ( .IN(n1851), .Q(g6258) );
  INVX1 U1729 ( .IN(n1891), .Q(n1909) );
  NOR2X1 U1730 ( .A(n1476), .B(n1511), .Q(n1557) );
  NAND2X1 U1731 ( .A(n1574), .B(n1575), .Q(n1472) );
  NOR2X1 U1732 ( .A(n1859), .B(n1482), .Q(n1571) );
  NOR2X1 U1733 ( .A(n1571), .B(n1482), .Q(n1483) );
  AND4X1 U1734 ( .A(n1548), .B(n1580), .C(n1849), .D(n1851), .Q(n1482)
         );
  AOI222X1 U1735 ( .A(n1485), .B(g1577), .C(n1482), .D(g296), .E(
        n1483), .F(g272), .Q(n1500) );
  AOI222X1 U1736 ( .A(n1485), .B(g1571), .C(n1482), .D(g290), .E(
        n1483), .F(g266), .Q(n1532) );
  NAND4X1 U1737 ( .A(n1551), .B(n1552), .C(n1553), .D(n1554), .Q(
        g10664) );
  INVX1 U1738 ( .IN(n1486), .Q(n577) );
  INVX1 U1739 ( .IN(n1909), .Q(n1854) );
  INVX1 U1740 ( .IN(n1909), .Q(n1853) );
  INVX1 U1741 ( .IN(n1565), .Q(n576) );
  NOR2X1 U1742 ( .A(n1566), .B(n1567), .Q(n1556) );
  INVX1 U1743 ( .IN(n1579), .Q(n572) );
  AND2X1 U1744 ( .A(n1574), .B(n1577), .Q(n1481) );
  NAND2X1 U1745 ( .A(n1547), .B(n1849), .Q(n1494) );
  INVX1 U1746 ( .IN(n1909), .Q(n1901) );
  INVX1 U1747 ( .IN(n1472), .Q(n580) );
  NAND4X1 U1748 ( .A(n1499), .B(n1500), .C(n1501), .D(n1502), .Q(
        g10722) );
  INVX1 U1749 ( .IN(n1909), .Q(n1902) );
  INVX1 U1750 ( .IN(n1895), .Q(n1921) );
  AND2X1 U1751 ( .A(n1574), .B(n1576), .Q(n1506) );
  INVX1 U1752 ( .IN(n1352), .Q(n1856) );
  AND2X1 U1753 ( .A(n1577), .B(n1544), .Q(n1476) );
  ISOLANDX1 U1754 ( .D(n1548), .ISO(n1545), .Q(n1479) );
  XOR3X1 U1755 ( .A(n1857), .B(n1243), .C(n1244), .Q(n1220) );
  XNOR3X1 U1756 ( .A(n1250), .B(n1251), .C(n1252), .Q(n1857) );
  XOR3X1 U1757 ( .A(n1858), .B(n1461), .C(n1462), .Q(n1459) );
  XNOR2X1 U1758 ( .A(g10722), .B(g10721), .Q(n1858) );
  NAND2X1 U1759 ( .A(n1971), .B(g10722), .Q(n1444) );
  INVX1 U1760 ( .IN(n1923), .Q(n1953) );
  INVX1 U1761 ( .IN(n1923), .Q(n1954) );
  INVX1 U1762 ( .IN(n1922), .Q(n1955) );
  INVX1 U1763 ( .IN(n1946), .Q(n1924) );
  INVX1 U1764 ( .IN(n1947), .Q(n1922) );
  INVX1 U1765 ( .IN(n1947), .Q(n1923) );
  INVX1 U1766 ( .IN(n1945), .Q(n1925) );
  INVX1 U1767 ( .IN(n1942), .Q(n1931) );
  INVX1 U1768 ( .IN(n1943), .Q(n1930) );
  INVX1 U1769 ( .IN(n1942), .Q(n1932) );
  INVX1 U1770 ( .IN(n1945), .Q(n1927) );
  INVX1 U1771 ( .IN(n1944), .Q(n1929) );
  INVX1 U1772 ( .IN(n1945), .Q(n1926) );
  INVX1 U1773 ( .IN(n1944), .Q(n1928) );
  INVX1 U1774 ( .IN(n1942), .Q(n1933) );
  INVX1 U1775 ( .IN(n1941), .Q(n1935) );
  INVX1 U1776 ( .IN(n1941), .Q(n1934) );
  INVX1 U1777 ( .IN(n1940), .Q(n1936) );
  INVX1 U1778 ( .IN(n1940), .Q(n1937) );
  INVX1 U1779 ( .IN(n1974), .Q(n1966) );
  INVX1 U1780 ( .IN(n1973), .Q(n1961) );
  INVX1 U1781 ( .IN(n1970), .Q(n1967) );
  INVX1 U1782 ( .IN(n1948), .Q(n1946) );
  INVX1 U1783 ( .IN(n1969), .Q(n1962) );
  INVX1 U1784 ( .IN(n1972), .Q(n1964) );
  INVX1 U1785 ( .IN(n1975), .Q(n1965) );
  INVX1 U1786 ( .IN(n1971), .Q(n1963) );
  INVX1 U1787 ( .IN(n1948), .Q(n1947) );
  INVX1 U1788 ( .IN(n1950), .Q(n1941) );
  INVX1 U1789 ( .IN(n1949), .Q(n1942) );
  INVX1 U1790 ( .IN(n1950), .Q(n1940) );
  INVX1 U1791 ( .IN(n1949), .Q(n1943) );
  INVX1 U1792 ( .IN(n1950), .Q(n1945) );
  INVX1 U1793 ( .IN(n1949), .Q(n1944) );
  INVX1 U1794 ( .IN(n1941), .Q(n1938) );
  INVX1 U1795 ( .IN(n1940), .Q(n1939) );
  INVX1 U1796 ( .IN(n1890), .Q(n1907) );
  INVX1 U1797 ( .IN(n1891), .Q(n1908) );
  ISOLANDX1 U1798 ( .D(n1567), .ISO(n1480), .Q(n1485) );
  NAND2X1 U1799 ( .A(n1557), .B(n1565), .Q(n1543) );
  INVX1 U1800 ( .IN(n1892), .Q(n1910) );
  INVX1 U1801 ( .IN(n1895), .Q(n1913) );
  INVX1 U1802 ( .IN(n1895), .Q(n1920) );
  INVX1 U1803 ( .IN(n1892), .Q(n1911) );
  INVX1 U1804 ( .IN(n1893), .Q(n1915) );
  INVX1 U1805 ( .IN(n1894), .Q(n1917) );
  INVX1 U1806 ( .IN(n1894), .Q(n1916) );
  INVX1 U1807 ( .IN(n1895), .Q(n1919) );
  INVX1 U1808 ( .IN(n1893), .Q(n1912) );
  INVX1 U1809 ( .IN(n1893), .Q(n1914) );
  INVX1 U1810 ( .IN(n1894), .Q(n1918) );
  INVX1 U1811 ( .IN(n1335), .Q(n522) );
  INVX1 U1812 ( .IN(n1982), .Q(n1971) );
  INVX1 U1813 ( .IN(n1981), .Q(n1972) );
  INVX1 U1814 ( .IN(n1980), .Q(n1973) );
  INVX1 U1815 ( .IN(n1982), .Q(n1970) );
  INVX1 U1816 ( .IN(n1979), .Q(n1974) );
  INVX1 U1817 ( .IN(n1952), .Q(n1948) );
  INVX1 U1818 ( .IN(n1983), .Q(n1969) );
  INVX1 U1819 ( .IN(n1979), .Q(n1975) );
  INVX1 U1820 ( .IN(n1978), .Q(n1976) );
  INVX1 U1821 ( .IN(n1951), .Q(n1950) );
  INVX1 U1822 ( .IN(n1951), .Q(n1949) );
  INVX1 U1823 ( .IN(n844), .Q(n605) );
  INVX1 U1824 ( .IN(n865), .Q(n597) );
  INVX1 U1825 ( .IN(n1959), .Q(n1880) );
  INVX1 U1826 ( .IN(n1959), .Q(g2355) );
  INVX1 U1827 ( .IN(n1144), .Q(n619) );
  INVX1 U1828 ( .IN(n1171), .Q(n553) );
  NOR4X1 U1829 ( .A(n1543), .B(n1491), .C(n1473), .D(n1512), .Q(n1509) );
  AND2X1 U1830 ( .A(n1576), .B(n1544), .Q(n1511) );
  AND2X1 U1831 ( .A(n1575), .B(n1548), .Q(n1480) );
  AO21X1 U1832 ( .A(n1576), .B(n1548), .C(n1480), .Q(n1567) );
  INVX1 U1833 ( .IN(n1889), .Q(n1905) );
  INVX1 U1834 ( .IN(n1899), .Q(n1890) );
  INVX1 U1835 ( .IN(n1444), .Q(n535) );
  NAND2X1 U1836 ( .A(n1902), .B(n625), .Q(n1360) );
  NAND2X1 U1837 ( .A(n1575), .B(n1544), .Q(n1565) );
  NAND2X1 U1838 ( .A(n524), .B(n617), .Q(n1335) );
  ISOLANDX1 U1839 ( .D(n1566), .ISO(n1479), .Q(n1486) );
  INVX1 U1840 ( .IN(n1896), .Q(n1894) );
  INVX1 U1841 ( .IN(n1897), .Q(n1895) );
  INVX1 U1842 ( .IN(n1897), .Q(n1893) );
  ISOLANDX1 U1843 ( .D(n1546), .ISO(n581), .Q(n1478) );
  INVX1 U1844 ( .IN(n1494), .Q(n579) );
  NOR2X1 U1845 ( .A(n1476), .B(n576), .Q(n1477) );
  INVX1 U1846 ( .IN(n1473), .Q(n573) );
  NAND2X1 U1847 ( .A(n1887), .B(n545), .Q(g10457) );
  NAND2X1 U1848 ( .A(n1886), .B(n544), .Q(g10455) );
  NAND2X1 U1849 ( .A(n1291), .B(n552), .Q(n1222) );
  NAND2X1 U1850 ( .A(n1887), .B(n546), .Q(g10459) );
  INVX1 U1851 ( .IN(n1988), .Q(n1968) );
  INVX1 U1852 ( .IN(n1984), .Q(n1982) );
  INVX1 U1853 ( .IN(n1985), .Q(n1981) );
  INVX1 U1854 ( .IN(n1985), .Q(n1980) );
  NAND2X1 U1855 ( .A(n1291), .B(n548), .Q(n1290) );
  INVX1 U1856 ( .IN(n1447), .Q(n532) );
  INVX1 U1857 ( .IN(n1445), .Q(n534) );
  NAND2X1 U1858 ( .A(n1887), .B(n548), .Q(g10465) );
  NAND2X1 U1859 ( .A(n1886), .B(n547), .Q(g10463) );
  NAND2X1 U1860 ( .A(n1886), .B(n552), .Q(g10377) );
  INVX1 U1861 ( .IN(n1983), .Q(n1977) );
  INVX1 U1862 ( .IN(n1986), .Q(n1978) );
  INVX1 U1863 ( .IN(n1986), .Q(n1979) );
  INVX1 U1864 ( .IN(n968), .Q(n1952) );
  NAND2X1 U1865 ( .A(n797), .B(n1395), .Q(n1291) );
  NAND2X1 U1866 ( .A(n1974), .B(n547), .Q(n1382) );
  INVX1 U1867 ( .IN(n1103), .Q(n557) );
  NAND2X1 U1868 ( .A(n668), .B(n649), .Q(n1101) );
  NAND2X1 U1869 ( .A(n623), .B(n715), .Q(n1144) );
  NAND2X1 U1870 ( .A(n715), .B(n598), .Q(n865) );
  NAND2X1 U1871 ( .A(n668), .B(n607), .Q(n844) );
  NAND2X1 U1872 ( .A(n555), .B(n1141), .Q(n1139) );
  NAND2X1 U1873 ( .A(n555), .B(n661), .Q(n1171) );
  INVX1 U1874 ( .IN(n1984), .Q(n1983) );
  INVX1 U1875 ( .IN(n968), .Q(n1951) );
  INVX1 U1876 ( .IN(n1592), .Q(n592) );
  ISOLANDX1 U1877 ( .D(n1137), .ISO(n1967), .Q(n1195) );
  NOR2X1 U1878 ( .A(n1026), .B(n649), .Q(n960) );
  NOR2X1 U1879 ( .A(n1641), .B(n1311), .Q(n1309) );
  INVX1 U1880 ( .IN(n866), .Q(n596) );
  INVX1 U1881 ( .IN(n845), .Q(n606) );
  INVX1 U1882 ( .IN(n850), .Q(n644) );
  INVX1 U1883 ( .IN(n855), .Q(n620) );
  INVX1 U1884 ( .IN(n1407), .Q(n662) );
  NOR2X1 U1885 ( .A(n529), .B(n1198), .Q(g5763) );
  NOR2X1 U1886 ( .A(n533), .B(n1181), .Q(g6392) );
  INVX1 U1887 ( .IN(n1005), .Q(n633) );
  INVX1 U1888 ( .IN(n1311), .Q(n611) );
  INVX1 U1889 ( .IN(n1295), .Q(n612) );
  INVX1 U1890 ( .IN(n830), .Q(n603) );
  INVX1 U1891 ( .IN(n875), .Q(n595) );
  INVX1 U1892 ( .IN(n933), .Q(n646) );
  INVX1 U1893 ( .IN(n863), .Q(n712) );
  INVX1 U1894 ( .IN(n908), .Q(n718) );
  AND3X1 U1895 ( .A(n1849), .B(n1851), .C(n1578), .Q(n1575) );
  NAND2X1 U1896 ( .A(n1581), .B(n1849), .Q(n1579) );
  NAND3X1 U1897 ( .A(n1579), .B(n1550), .C(n1556), .Q(n1473) );
  AND3X1 U1898 ( .A(n1831), .B(n1841), .C(n842), .Q(n1395) );
  AND4X1 U1899 ( .A(n1571), .B(n583), .C(n1572), .D(n1573), .Q(n1546)
         );
  NOR2X1 U1900 ( .A(n1507), .B(n1530), .Q(n1572) );
  NOR4X1 U1901 ( .A(n1481), .B(n1506), .C(n580), .D(n1508), .Q(n1573)
         );
  INVX1 U1902 ( .IN(n1239), .Q(n1899) );
  INVX1 U1903 ( .IN(n1900), .Q(n1889) );
  INVX1 U1904 ( .IN(n1239), .Q(n1900) );
  AO21X1 U1905 ( .A(n1577), .B(n1548), .C(n1479), .Q(n1566) );
  XOR3X1 U1906 ( .A(n1245), .B(n1246), .C(n1247), .Q(n1243) );
  XOR2X1 U1907 ( .A(n1253), .B(n1254), .Q(n1251) );
  ISOLANDX1 U1908 ( .D(n1544), .ISO(n1545), .Q(n1512) );
  ISOLANDX1 U1909 ( .D(n1574), .ISO(n1545), .Q(n1530) );
  AND3X1 U1910 ( .A(n1548), .B(n1580), .C(n1396), .Q(n1859) );
  NAND4X1 U1911 ( .A(n1546), .B(n1495), .C(n1494), .D(n1541), .Q(
        n1491) );
  AND2X1 U1912 ( .A(n1396), .B(n1578), .Q(n1576) );
  XOR2X1 U1913 ( .A(n1248), .B(n1249), .Q(n1246) );
  NAND4X1 U1914 ( .A(n1444), .B(n1445), .C(n1446), .D(n1447), .Q(
        n1440) );
  NAND2X1 U1915 ( .A(n1972), .B(n1448), .Q(n1446) );
  NAND4X1 U1916 ( .A(n547), .B(n545), .C(n548), .D(n1449), .Q(n1448)
         );
  NOR2X1 U1917 ( .A(g10663), .B(g10664), .Q(n1449) );
  XOR2X1 U1918 ( .A(n793), .B(n794), .Q(g11163) );
  OA21X1 U1919 ( .A(n1302), .B(n1606), .C(n1903), .Q(n1349) );
  INVX1 U1920 ( .IN(n1239), .Q(n1898) );
  INVX1 U1921 ( .IN(n1239), .Q(n1897) );
  INVX1 U1922 ( .IN(n1239), .Q(n1896) );
  NOR2X1 U1923 ( .A(n1344), .B(n1345), .Q(g11380) );
  OA21X1 U1924 ( .A(n1302), .B(n527), .C(n1606), .Q(n1344) );
  NOR2X1 U1925 ( .A(n1348), .B(n1345), .Q(g11372) );
  OA221X1 U1926 ( .A(n1349), .B(n1594), .C(n527), .D(n1350), .E(
        n1306), .Q(n1348) );
  NAND2X1 U1927 ( .A(n1884), .B(n1594), .Q(n1350) );
  XOR2X1 U1928 ( .A(n544), .B(n545), .Q(n1461) );
  XOR3X1 U1929 ( .A(n1463), .B(n548), .C(g10664), .Q(n1462) );
  NOR2X1 U1930 ( .A(n1353), .B(n1345), .Q(g11340) );
  XOR2X1 U1931 ( .A(n527), .B(n1884), .Q(n1353) );
  INVX1 U1932 ( .IN(n1464), .Q(g10628) );
  INVX1 U1933 ( .IN(n1541), .Q(n581) );
  NAND4X1 U1934 ( .A(n1556), .B(n1478), .C(n1557), .D(n1550), .Q(
        n1552) );
  INVX1 U1935 ( .IN(n1550), .Q(n575) );
  INVX1 U1936 ( .IN(n1495), .Q(n578) );
  INVX1 U1937 ( .IN(n793), .Q(n542) );
  NAND2X1 U1938 ( .A(n1974), .B(g10664), .Q(n1455) );
  AO221X1 U1939 ( .A(n1371), .B(g10726), .C(n1372), .D(g10664), .E(
        n1653), .Q(n1369) );
  AO221X1 U1940 ( .A(n1373), .B(g10720), .C(n1374), .D(g10722), .E(
        n1653), .Q(n1367) );
  AO22X1 U1941 ( .A(n662), .B(n1069), .C(n1454), .D(n1407), .Q(n1452)
         );
  NAND2X1 U1942 ( .A(n1611), .B(n1455), .Q(n1454) );
  AO22X1 U1943 ( .A(n662), .B(n1075), .C(n1404), .D(n535), .Q(n1405)
         );
  INVX1 U1944 ( .IN(g10720), .Q(n545) );
  NAND2X1 U1945 ( .A(n1973), .B(g10721), .Q(n1447) );
  NAND2X1 U1946 ( .A(n1968), .B(g10719), .Q(n1445) );
  INVX1 U1947 ( .IN(g10724), .Q(n547) );
  INVX1 U1948 ( .IN(g10719), .Q(n544) );
  INVX1 U1949 ( .IN(g10726), .Q(n548) );
  NAND2X1 U1950 ( .A(n1969), .B(g10720), .Q(n1414) );
  INVX1 U1951 ( .IN(n1987), .Q(n1984) );
  INVX1 U1952 ( .IN(n1987), .Q(n1985) );
  AO22X1 U1953 ( .A(n662), .B(n1067), .C(n1404), .D(n532), .Q(n1408)
         );
  AO22X1 U1954 ( .A(n662), .B(n1063), .C(n1418), .D(n1407), .Q(n1410)
         );
  NAND2X1 U1955 ( .A(n1416), .B(n545), .Q(n1418) );
  AO22X1 U1956 ( .A(n662), .B(n1084), .C(n1404), .D(n534), .Q(n1412)
         );
  AO22X1 U1957 ( .A(n662), .B(n1077), .C(n1415), .D(n1407), .Q(n1411)
         );
  NAND2X1 U1958 ( .A(n1416), .B(n544), .Q(n1415) );
  INVX1 U1959 ( .IN(g10663), .Q(n552) );
  INVX1 U1960 ( .IN(g10721), .Q(n546) );
  INVX1 U1961 ( .IN(n1255), .Q(n549) );
  AO22X1 U1962 ( .A(n662), .B(n1082), .C(n1413), .D(n1407), .Q(n1409)
         );
  NAND2X1 U1963 ( .A(n1611), .B(n1414), .Q(n1413) );
  XOR2X1 U1964 ( .A(g10724), .B(g10663), .Q(n1463) );
  NAND2X1 U1965 ( .A(n550), .B(n1229), .Q(n1225) );
  NAND2X1 U1966 ( .A(n1261), .B(n1262), .Q(n1259) );
  INVX1 U1967 ( .IN(n1227), .Q(n550) );
  NOR2X1 U1968 ( .A(n1965), .B(n1113), .Q(n1120) );
  INVX1 U1969 ( .IN(n1867), .Q(n1887) );
  INVX1 U1970 ( .IN(n1867), .Q(n1886) );
  NAND2X1 U1971 ( .A(n1113), .B(n1114), .Q(n1103) );
  AND4X1 U1972 ( .A(n1396), .B(n1847), .C(n1845), .D(n1843), .Q(n797)
         );
  INVX1 U1973 ( .IN(n1988), .Q(n1986) );
  AO221X1 U1974 ( .A(n1404), .B(g10663), .C(n662), .D(n1088), .E(
        n1450), .Q(n1453) );
  AO22X1 U1975 ( .A(n662), .B(n1080), .C(n1404), .D(n1382), .Q(n1402)
         );
  AO221X1 U1976 ( .A(n1404), .B(g10726), .C(n662), .D(n1086), .E(
        n1450), .Q(n1417) );
  NOR2X1 U1977 ( .A(n1217), .B(n1961), .Q(g5392) );
  NOR2X1 U1978 ( .A(n1683), .B(n1961), .Q(n1198) );
  NOR2X1 U1979 ( .A(n594), .B(n1961), .Q(n1181) );
  NOR2X1 U1980 ( .A(n1362), .B(n1363), .Q(n1352) );
  NAND2X1 U1981 ( .A(n560), .B(n744), .Q(n968) );
  INVX1 U1982 ( .IN(n1059), .Q(n533) );
  INVX1 U1983 ( .IN(n1236), .Q(n529) );
  NAND4X1 U1984 ( .A(n844), .B(n805), .C(n952), .D(n953), .Q(n845) );
  NOR2X1 U1985 ( .A(n954), .B(n720), .Q(n952) );
  NAND4X1 U1986 ( .A(n865), .B(n815), .C(n916), .D(n715), .Q(n866) );
  ISOLANDX1 U1987 ( .D(n822), .ISO(n809), .Q(n916) );
  NAND4X1 U1988 ( .A(n1684), .B(n1623), .C(n1601), .D(n1590), .Q(
        n1289) );
  NAND2X1 U1989 ( .A(n648), .B(n958), .Q(n850) );
  NAND2X1 U1990 ( .A(n622), .B(n918), .Q(n855) );
  NAND3X1 U1991 ( .A(n1833), .B(n1775), .C(n842), .Q(g9961) );
  NOR2X1 U1992 ( .A(n891), .B(n1657), .Q(n875) );
  NOR2X1 U1993 ( .A(n949), .B(n1656), .Q(n933) );
  NOR2X1 U1994 ( .A(n1054), .B(n1117), .Q(n1116) );
  NOR2X1 U1995 ( .A(n607), .B(n805), .Q(n830) );
  NAND2X1 U1996 ( .A(n1648), .B(n1611), .Q(n1407) );
  NOR2X1 U1997 ( .A(n650), .B(n954), .Q(n1035) );
  NOR2X1 U1998 ( .A(n624), .B(n1032), .Q(n1039) );
  NAND2X1 U1999 ( .A(n675), .B(n1594), .Q(n1311) );
  NAND2X1 U2000 ( .A(n985), .B(n1658), .Q(n1005) );
  NAND2X1 U2001 ( .A(n674), .B(n1594), .Q(n1295) );
  NAND2X1 U2002 ( .A(n1773), .B(n1665), .Q(g8352) );
  NAND2X1 U2003 ( .A(n1773), .B(n1669), .Q(g8349) );
  NAND2X1 U2004 ( .A(n1773), .B(n1666), .Q(g8335) );
  NAND2X1 U2005 ( .A(n1773), .B(n1664), .Q(g8328) );
  NAND2X1 U2006 ( .A(n1773), .B(n1667), .Q(g8318) );
  NAND2X1 U2007 ( .A(n1773), .B(n1668), .Q(g8313) );
  NAND2X1 U2008 ( .A(n1773), .B(n1671), .Q(g8347) );
  NAND2X1 U2009 ( .A(n1773), .B(n1670), .Q(g8340) );
  NAND2X1 U2010 ( .A(n1773), .B(n1672), .Q(g8331) );
  NAND2X1 U2011 ( .A(n1773), .B(n1673), .Q(g8323) );
  NAND2X1 U2012 ( .A(n1773), .B(n1674), .Q(g8316) );
  NAND3X1 U2013 ( .A(n814), .B(n815), .C(n826), .Q(n863) );
  NAND3X1 U2014 ( .A(n831), .B(n832), .C(n966), .Q(n908) );
  NOR2X1 U2015 ( .A(n1029), .B(n1622), .Q(n1191) );
  NOR2X1 U2016 ( .A(n1593), .B(n1607), .Q(n834) );
  NOR2X1 U2017 ( .A(n1634), .B(n1957), .Q(n1137) );
  INVX1 U2018 ( .IN(n1169), .Q(n538) );
  INVX1 U2019 ( .IN(n1167), .Q(n539) );
  NOR2X1 U2020 ( .A(n1963), .B(n1159), .Q(n1173) );
  NAND4X1 U2021 ( .A(n721), .B(n1593), .C(n1609), .D(n1645), .Q(n1026) );
  NAND4X1 U2022 ( .A(n648), .B(n718), .C(n1615), .D(n1662), .Q(n950)
         );
  NAND4X1 U2023 ( .A(n622), .B(n712), .C(n1616), .D(n1663), .Q(n892)
         );
  OA221X1 U2024 ( .A(n599), .B(n810), .C(n811), .D(n1605), .E(n1880), 
        .Q(g9272) );
  NAND2X1 U2025 ( .A(n715), .B(n1605), .Q(n810) );
  INVX1 U2026 ( .IN(n811), .Q(n599) );
  NAND2X1 U2027 ( .A(n812), .B(n813), .Q(n811) );
  NOR2X1 U2028 ( .A(n1659), .B(n1172), .Q(n1141) );
  NOR2X1 U2029 ( .A(n1183), .B(n1714), .Q(g6179) );
  INVX1 U2030 ( .IN(n1142), .Q(n517) );
  ISOLANDX1 U2031 ( .D(n1057), .ISO(n1054), .Q(n1056) );
  NOR2X1 U2032 ( .A(n1626), .B(n1117), .Q(n1057) );
  INVX1 U2033 ( .IN(n899), .Q(n648) );
  INVX1 U2034 ( .IN(n853), .Q(n622) );
  ISOLANDX1 U2035 ( .D(n1404), .ISO(n1969), .Q(n1450) );
  OR2X1 U2036 ( .A(n1616), .B(n922), .Q(n925) );
  OR2X1 U2037 ( .A(n1615), .B(n846), .Q(n849) );
  NOR2X1 U2038 ( .A(n1306), .B(n1307), .Q(n1304) );
  NOR3X1 U2039 ( .A(n598), .B(n1605), .C(n826), .Q(n820) );
  NOR2X1 U2040 ( .A(n1264), .B(n1263), .Q(n1258) );
  AO21X1 U2041 ( .A(n605), .B(n951), .C(n606), .Q(g8883) );
  XOR2X1 U2042 ( .A(n1656), .B(n955), .Q(n951) );
  NAND2X1 U2043 ( .A(n850), .B(n956), .Q(n955) );
  NAND3X1 U2044 ( .A(n950), .B(n949), .C(n957), .Q(n956) );
  AO21X1 U2045 ( .A(n597), .B(n893), .C(n596), .Q(g8937) );
  XOR2X1 U2046 ( .A(n1657), .B(n894), .Q(n893) );
  NAND2X1 U2047 ( .A(n855), .B(n895), .Q(n894) );
  NAND3X1 U2048 ( .A(n892), .B(n891), .C(n896), .Q(n895) );
  AO21X1 U2049 ( .A(n597), .B(n887), .C(n596), .Q(g8938) );
  XOR2X1 U2050 ( .A(n1675), .B(n888), .Q(n887) );
  NAND2X1 U2051 ( .A(n855), .B(n889), .Q(n888) );
  NAND3X1 U2052 ( .A(n600), .B(n595), .C(n890), .Q(n889) );
  AO21X1 U2053 ( .A(n605), .B(n945), .C(n606), .Q(g8885) );
  XOR2X1 U2054 ( .A(n1676), .B(n946), .Q(n945) );
  NAND2X1 U2055 ( .A(n850), .B(n947), .Q(n946) );
  NAND3X1 U2056 ( .A(n645), .B(n646), .C(n948), .Q(n947) );
  INVX1 U2057 ( .IN(n1054), .Q(n555) );
  NAND3X1 U2058 ( .A(n814), .B(n815), .C(n816), .Q(n813) );
  OR2X1 U2059 ( .A(n817), .B(n1643), .Q(n816) );
  NBUFFX1 U2060 ( .IN(n1960), .Q(n1957) );
  NOR2X1 U2061 ( .A(n1884), .B(n1311), .Q(n1313) );
  NBUFFX1 U2062 ( .IN(n1960), .Q(n1958) );
  NOR2X1 U2063 ( .A(n1038), .B(n623), .Q(n929) );
  NAND2X1 U2064 ( .A(n1593), .B(n1644), .Q(n964) );
  NAND2X1 U2065 ( .A(n1263), .B(n1264), .Q(n1262) );
  NOR2X1 U2066 ( .A(n1965), .B(n1596), .Q(g4506) );
  NOR2X1 U2067 ( .A(n1964), .B(n1602), .Q(g6193) );
  NOR2X1 U2068 ( .A(n1964), .B(n1619), .Q(g6331) );
  NOR2X1 U2069 ( .A(n1965), .B(n1660), .Q(g4490) );
  NOR2X1 U2070 ( .A(n1965), .B(n1618), .Q(g4471) );
  NOR2X1 U2071 ( .A(n1964), .B(n1700), .Q(g6332) );
  NOR2X1 U2072 ( .A(n1964), .B(n1617), .Q(g4498) );
  NOR2X1 U2073 ( .A(n1965), .B(n1708), .Q(g4473) );
  NOR2X1 U2074 ( .A(n1964), .B(n1685), .Q(g4342) );
  NOR2X1 U2075 ( .A(n1964), .B(n1705), .Q(g4477) );
  NOR2X1 U2076 ( .A(n1965), .B(n1597), .Q(g4484) );
  NOR2X1 U2077 ( .A(n1963), .B(n1624), .Q(g6828) );
  NOR2X1 U2078 ( .A(n1964), .B(n1627), .Q(g6205) );
  NOR2X1 U2079 ( .A(n1962), .B(n1073), .Q(g8047) );
  XOR2X1 U2080 ( .A(n1704), .B(g6035), .Q(n1073) );
  NOR2X1 U2081 ( .A(n1962), .B(n1081), .Q(g8042) );
  XOR2X1 U2082 ( .A(n1703), .B(n1082), .Q(n1081) );
  NOR2X1 U2083 ( .A(n1963), .B(n1625), .Q(g6820) );
  NOR2X1 U2084 ( .A(n1963), .B(n1603), .Q(g6334) );
  NOR2X1 U2085 ( .A(n1965), .B(n1661), .Q(g4465) );
  NOR2X1 U2086 ( .A(n1963), .B(n1688), .Q(g6834) );
  NOR2X1 U2087 ( .A(n1963), .B(n1598), .Q(g6840) );
  NOR2X1 U2088 ( .A(n1964), .B(n1628), .Q(g6180) );
  NOR2X1 U2089 ( .A(n1965), .B(n1706), .Q(g4480) );
  NOR2X1 U2090 ( .A(n1964), .B(n1710), .Q(g6224) );
  NOR2X1 U2091 ( .A(n1963), .B(n1711), .Q(g6839) );
  NOR2X1 U2092 ( .A(n1964), .B(n1678), .Q(g6333) );
  NOR2X1 U2093 ( .A(n1963), .B(n1629), .Q(g6841) );
  NOR2X1 U2094 ( .A(n1965), .B(n1686), .Q(g4340) );
  NOR2X1 U2095 ( .A(n1963), .B(n1687), .Q(g6830) );
  NOR2X1 U2096 ( .A(n1953), .B(n1648), .Q(g4500) );
  NOR2X1 U2097 ( .A(n1654), .B(n1216), .Q(g5390) );
  NOR2X1 U2098 ( .A(n1614), .B(n1216), .Q(g5148) );
  NOR2X1 U2099 ( .A(n1677), .B(n1216), .Q(g5173) );
  NOR2X1 U2100 ( .A(n1658), .B(n1216), .Q(g5126) );
  NOR2X1 U2101 ( .A(n1630), .B(n1040), .Q(g8254) );
  NOR2X1 U2102 ( .A(n1604), .B(n1040), .Q(g8147) );
  NOR2X1 U2103 ( .A(n1591), .B(n1040), .Q(g8250) );
  NOR2X1 U2104 ( .A(n1712), .B(n1040), .Q(g8260) );
  NOR2X1 U2105 ( .A(n644), .B(n912), .Q(n911) );
  NOR2X1 U2106 ( .A(n620), .B(n869), .Q(n868) );
  NBUFFX1 U2107 ( .IN(n1960), .Q(n1959) );
  NAND2X1 U2108 ( .A(n830), .B(n1713), .Q(n803) );
  NAND2X1 U2109 ( .A(n685), .B(n1595), .Q(n1128) );
  INVX1 U2110 ( .IN(n1183), .Q(n519) );
  NOR3X1 U2111 ( .A(n1953), .B(g4089), .C(n561), .Q(g5083) );
  NOR2X1 U2112 ( .A(n1885), .B(n1170), .Q(g6516) );
  OA22X1 U2113 ( .A(n1141), .B(n1171), .C(n554), .D(n1659), .Q(n1170)
         );
  INVX1 U2114 ( .IN(n1139), .Q(n554) );
  NOR2X1 U2115 ( .A(n1885), .B(n1115), .Q(g7541) );
  OA22X1 U2116 ( .A(n1057), .B(n556), .C(n1056), .D(n1626), .Q(n1115)
         );
  INVX1 U2117 ( .IN(n1116), .Q(n556) );
  NAND2X1 U2118 ( .A(n1605), .B(n1643), .Q(n928) );
  NOR2X1 U2119 ( .A(n1957), .B(n839), .Q(g9110) );
  XOR2X1 U2120 ( .A(n1607), .B(n840), .Q(n839) );
  NAND3X1 U2121 ( .A(n837), .B(n603), .C(n841), .Q(n840) );
  NAND2X1 U2122 ( .A(n804), .B(n719), .Q(n841) );
  INVX1 U2123 ( .IN(n1160), .Q(n667) );
  INVX1 U2124 ( .IN(n1148), .Q(n711) );
  NAND2X1 U2125 ( .A(n1160), .B(n1701), .Q(g6672) );
  NAND2X1 U2126 ( .A(n795), .B(n796), .Q(n1585) );
  NAND2X1 U2127 ( .A(n797), .B(n798), .Q(n1587) );
  NAND2X1 U2128 ( .A(n795), .B(n798), .Q(n1588) );
  NAND2X1 U2129 ( .A(n797), .B(n796), .Q(n1586) );
  INVX1 U2130 ( .IN(n1016), .Q(n650) );
  INVX1 U2131 ( .IN(n1031), .Q(n624) );
  NAND4X1 U2132 ( .A(n1380), .B(n822), .C(n1038), .D(n920), .Q(n1379)
         );
  NAND2X1 U2133 ( .A(n713), .B(n1605), .Q(n814) );
  NAND2X1 U2134 ( .A(n719), .B(n1593), .Q(n831) );
  INVX1 U2135 ( .IN(n1046), .Q(n537) );
  INVX1 U2136 ( .IN(n1025), .Q(n719) );
  INVX1 U2137 ( .IN(n1306), .Q(n610) );
  INVX1 U2138 ( .IN(n978), .Q(n631) );
  INVX1 U2139 ( .IN(n954), .Q(n668) );
  INVX1 U2140 ( .IN(n1109), .Q(n540) );
  INVX1 U2141 ( .IN(n1032), .Q(n715) );
  INVX1 U2142 ( .IN(n1325), .Q(n674) );
  INVX1 U2143 ( .IN(n1307), .Q(n675) );
  INVX1 U2144 ( .IN(n920), .Q(n713) );
  INVX1 U2145 ( .IN(n877), .Q(n600) );
  INVX1 U2146 ( .IN(n935), .Q(n645) );
  INVX1 U2147 ( .IN(n1092), .Q(n630) );
  INVX1 U2148 ( .IN(n953), .Q(n717) );
  OAI21X1 U2149 ( .A(n915), .B(n865), .C(n866), .Q(g8921) );
  OA22X1 U2150 ( .A(n922), .B(n923), .C(n924), .D(n1616), .Q(n915) );
  NAND2X1 U2151 ( .A(n855), .B(n925), .Q(n923) );
  NOR2X1 U2152 ( .A(n620), .B(n925), .Q(n924) );
  OAI21X1 U2153 ( .A(n843), .B(n844), .C(n845), .Q(g8973) );
  OA22X1 U2154 ( .A(n846), .B(n847), .C(n848), .D(n1615), .Q(n843) );
  NAND2X1 U2155 ( .A(n850), .B(n849), .Q(n847) );
  NOR2X1 U2156 ( .A(n644), .B(n849), .Q(n848) );
  OAI21X1 U2157 ( .A(n909), .B(n844), .C(n845), .Q(g8922) );
  OA22X1 U2158 ( .A(n647), .B(n910), .C(n911), .D(n1662), .Q(n909) );
  INVX1 U2159 ( .IN(n913), .Q(n647) );
  NAND2X1 U2160 ( .A(n850), .B(n912), .Q(n910) );
  OAI21X1 U2161 ( .A(n864), .B(n865), .C(n866), .Q(g8943) );
  OA22X1 U2162 ( .A(n621), .B(n867), .C(n868), .D(n1663), .Q(n864) );
  INVX1 U2163 ( .IN(n870), .Q(n621) );
  NAND2X1 U2164 ( .A(n855), .B(n869), .Q(n867) );
  INVX1 U2165 ( .IN(n1384), .Q(n536) );
  INVX1 U2166 ( .IN(n1042), .Q(n520) );
  INVX1 U2167 ( .IN(n1119), .Q(n685) );
  OA221X1 U2168 ( .A(n604), .B(n827), .C(n828), .D(n1593), .E(g2355), 
        .Q(g9150) );
  NAND2X1 U2169 ( .A(n668), .B(n1593), .Q(n827) );
  INVX1 U2170 ( .IN(n828), .Q(n604) );
  OA21X1 U2171 ( .A(n607), .B(n829), .C(n803), .Q(n828) );
  INVX1 U2172 ( .IN(n966), .Q(n721) );
  INVX1 U2173 ( .IN(n959), .Q(n649) );
  INVX1 U2174 ( .IN(n993), .Q(n632) );
  INVX1 U2175 ( .IN(n1318), .Q(n609) );
  INVX1 U2176 ( .IN(n999), .Q(n634) );
  INVX1 U2177 ( .IN(n926), .Q(n623) );
  INVX1 U2178 ( .IN(n832), .Q(n720) );
  INVX1 U2179 ( .IN(n1302), .Q(n614) );
  INVX1 U2180 ( .IN(n804), .Q(n607) );
  INVX1 U2181 ( .IN(n812), .Q(n598) );
  INVX1 U2182 ( .IN(n1114), .Q(n629) );
  INVX1 U2183 ( .IN(n1110), .Q(n665) );
  INVX1 U2184 ( .IN(n974), .Q(n564) );
  INVX1 U2185 ( .IN(n995), .Q(n568) );
  INVX1 U2186 ( .IN(n1001), .Q(n566) );
  INVX1 U2187 ( .IN(n981), .Q(n563) );
  INVX1 U2188 ( .IN(n989), .Q(n567) );
  INVX1 U2189 ( .IN(n1007), .Q(n569) );
  INVX1 U2190 ( .IN(n1012), .Q(n565) );
  INVX1 U2191 ( .IN(n1420), .Q(n625) );
  INVX1 U2192 ( .IN(n1166), .Q(n518) );
  INVX1 U2193 ( .IN(n1875), .Q(n1888) );
  NOR2X1 U2194 ( .A(n1126), .B(n1101), .Q(g7137) );
  OA22X1 U2195 ( .A(n1127), .B(n1709), .C(n651), .D(n1128), .Q(n1126)
         );
  INVX1 U2196 ( .IN(n1129), .Q(n651) );
  NOR2X1 U2197 ( .A(n1701), .B(n1129), .Q(n1127) );
  NOR2X1 U2198 ( .A(n1130), .B(n1101), .Q(g7134) );
  OA21X1 U2199 ( .A(n685), .B(n1595), .C(n1128), .Q(n1130) );
  INVX1 U2200 ( .IN(n1217), .Q(n725) );
  NOR4X1 U2201 ( .A(n1712), .B(n1630), .C(n1604), .D(n1591), .Q(g3381) );
  NOR2X1 U2202 ( .A(n592), .B(n1664), .Q(g6638) );
  NOR2X1 U2203 ( .A(n592), .B(n1665), .Q(g6531) );
  NOR2X1 U2204 ( .A(n592), .B(n1666), .Q(g6653) );
  NOR2X1 U2205 ( .A(n592), .B(n1667), .Q(g6627) );
  NOR2X1 U2206 ( .A(n592), .B(n1668), .Q(g6621) );
  NOR2X1 U2207 ( .A(n592), .B(n1669), .Q(g6526) );
  NAND2X1 U2208 ( .A(n1148), .B(n1642), .Q(g6755) );
  NOR2X1 U2209 ( .A(n555), .B(n1601), .Q(g10780) );
  NOR2X1 U2210 ( .A(n555), .B(n1623), .Q(g10785) );
  NOR2X1 U2211 ( .A(n555), .B(n1684), .Q(g10784) );
  NOR2X1 U2212 ( .A(n555), .B(n1590), .Q(g10782) );
  INVX1 U2213 ( .IN(n1451), .Q(n561) );
  NAND2X1 U2214 ( .A(n1670), .B(n1592), .Q(g7219) );
  NAND2X1 U2215 ( .A(n1671), .B(n1592), .Q(g7143) );
  NAND2X1 U2216 ( .A(n1672), .B(n1592), .Q(g7204) );
  NAND2X1 U2217 ( .A(n1673), .B(n1592), .Q(g7189) );
  NAND2X1 U2218 ( .A(n1674), .B(n1592), .Q(g7183) );
  INVX1 U2219 ( .IN(n1228), .Q(n687) );
  INVX1 U2220 ( .IN(n1338), .Q(n616) );
  INVX1 U2221 ( .IN(n1342), .Q(n617) );
  INVX1 U2222 ( .IN(n1172), .Q(n661) );
  OA22X1 U2223 ( .A(n577), .B(n1632), .C(n583), .D(DFF_228_n1), .Q(
        n1499) );
  AOI221X1 U2224 ( .A(n1479), .B(g1558), .C(n1480), .D(g1601), .E(
        n1513), .Q(n1501) );
  NAND2X1 U2225 ( .A(g6257), .B(n1581), .Q(n1550) );
  NOR3X1 U2226 ( .A(g833), .B(g841), .C(g837), .Q(n1441) );
  NOR4X1 U2227 ( .A(n1443), .B(g853), .C(g861), .D(g857), .Q(n1442)
         );
  NAND2X1 U2228 ( .A(g6263), .B(n1775), .Q(n1484) );
  NAND2X1 U2229 ( .A(n1547), .B(g6257), .Q(n1495) );
  NOR2X1 U2230 ( .A(n1849), .B(g6258), .Q(n1396) );
  NOR2X1 U2231 ( .A(g6263), .B(g6256), .Q(n1583) );
  NOR2X1 U2232 ( .A(n1847), .B(g6260), .Q(n1580) );
  AND4X1 U2233 ( .A(n1548), .B(g6258), .C(n1847), .D(n1845), .Q(n1547)
         );
  AND3X1 U2234 ( .A(n842), .B(n1831), .C(g6262), .Q(n796) );
  AND3X1 U2235 ( .A(n842), .B(n1841), .C(g6261), .Q(n798) );
  NOR2X1 U2236 ( .A(n1845), .B(g6259), .Q(n1578) );
  NOR2X1 U2237 ( .A(n1843), .B(g6256), .Q(n1569) );
  AND3X1 U2238 ( .A(g6257), .B(g6258), .C(n1580), .Q(n1577) );
  AO222X1 U2239 ( .A(n572), .B(g1753), .C(n579), .D(n1631), .E(n575), 
        .F(g1730), .Q(n1513) );
  AO21X1 U2240 ( .A(g318), .B(n1905), .C(n1315), .Q(n1247) );
  OA221X1 U2241 ( .A(n1316), .B(g486), .C(n1621), .D(n1317), .E(
        n1902), .Q(n1315) );
  NAND2X1 U2242 ( .A(n609), .B(n1883), .Q(n1317) );
  NOR2X1 U2243 ( .A(n1641), .B(n1318), .Q(n1316) );
  AO21X1 U2244 ( .A(g330), .B(n1904), .C(n1299), .Q(n1252) );
  OA221X1 U2245 ( .A(n1300), .B(g506), .C(n1600), .D(n1301), .E(
        n1854), .Q(n1299) );
  NAND2X1 U2246 ( .A(n614), .B(n1606), .Q(n1301) );
  NOR2X1 U2247 ( .A(g471), .B(n1302), .Q(n1300) );
  AO22X1 U2248 ( .A(n1592), .B(g336), .C(n1219), .D(n592), .Q(g11647)
         );
  OAI22X1 U2249 ( .A(n551), .B(n1220), .C(n1221), .D(n1222), .Q(n1219) );
  INVX1 U2250 ( .IN(n1222), .Q(n551) );
  AO22X1 U2251 ( .A(g345), .B(n1592), .C(n1237), .D(n592), .Q(g11625)
         );
  XOR2X1 U2252 ( .A(n1220), .B(n1221), .Q(n1237) );
  AO21X1 U2253 ( .A(g324), .B(n1906), .C(n1308), .Q(n1249) );
  OA221X1 U2254 ( .A(n1309), .B(g496), .C(n1689), .D(n1310), .E(
        n1901), .Q(n1308) );
  NAND2X1 U2255 ( .A(n611), .B(n1884), .Q(n1310) );
  AO21X1 U2256 ( .A(g309), .B(n1904), .C(n1292), .Q(n1254) );
  OA221X1 U2257 ( .A(n1293), .B(g516), .C(n1620), .D(n1294), .E(
        n1901), .Q(n1292) );
  NAND2X1 U2258 ( .A(n1884), .B(n612), .Q(n1294) );
  NOR2X1 U2259 ( .A(n1295), .B(n1641), .Q(n1293) );
  AO21X1 U2260 ( .A(g315), .B(n1907), .C(n1319), .Q(n1245) );
  OA221X1 U2261 ( .A(n1320), .B(g481), .C(n1680), .D(n1321), .E(
        n1901), .Q(n1319) );
  NAND2X1 U2262 ( .A(n609), .B(n1641), .Q(n1321) );
  NOR2X1 U2263 ( .A(n1884), .B(n1318), .Q(n1320) );
  AO21X1 U2264 ( .A(g327), .B(n1905), .C(n1303), .Q(n1250) );
  OA221X1 U2265 ( .A(n1304), .B(g501), .C(n1690), .D(n1305), .E(
        n1901), .Q(n1303) );
  NAND2X1 U2266 ( .A(n675), .B(n610), .Q(n1305) );
  AO21X1 U2267 ( .A(g321), .B(n1908), .C(n1312), .Q(n1248) );
  OA221X1 U2268 ( .A(n1313), .B(g491), .C(n1691), .D(n1314), .E(
        n1901), .Q(n1312) );
  NAND2X1 U2269 ( .A(n611), .B(n1641), .Q(n1314) );
  AO21X1 U2270 ( .A(g333), .B(n1906), .C(n1296), .Q(n1253) );
  OA221X1 U2271 ( .A(n1297), .B(g511), .C(n1679), .D(n1298), .E(
        n1901), .Q(n1296) );
  NAND2X1 U2272 ( .A(n612), .B(n1641), .Q(n1298) );
  NOR2X1 U2273 ( .A(n1884), .B(n1295), .Q(n1297) );
  NOR3X1 U2274 ( .A(n1503), .B(n1504), .C(n1505), .Q(n1502) );
  AO222X1 U2275 ( .A(g986), .B(n1506), .C(g959), .D(n580), .E(g4199), 
        .F(n1481), .Q(n1505) );
  AOI22X1 U2276 ( .A(n1506), .B(g947), .C(n1483), .D(g284), .Q(n1553)
         );
  OA221X1 U2277 ( .A(n583), .B(DFF_319_n1), .C(n1550), .D(n1633), 
        .E(n1555), .Q(n1554) );
  NOR2X1 U2278 ( .A(n1545), .B(n1831), .Q(n1570) );
  AOI22X1 U2279 ( .A(n1860), .B(n1861), .C(n1861), .D(n1459), .Q(n793) );
  OR2X1 U2280 ( .A(g32), .B(n583), .Q(n1860) );
  OAI21X1 U2281 ( .A(g32), .B(n583), .C(n1459), .Q(n1861) );
  AO221X1 U2282 ( .A(g5392), .B(g10663), .C(n535), .D(n1198), .E(
        n1465), .Q(n794) );
  AO222X1 U2283 ( .A(n1466), .B(n1977), .C(g2648), .D(n530), .E(n529), .F(g10724), .Q(n1465) );
  NOR2X1 U2284 ( .A(g105), .B(n548), .Q(n1466) );
  INVX1 U2285 ( .IN(n1455), .Q(n530) );
  NAND3X1 U2286 ( .A(n1853), .B(n1419), .C(n1420), .Q(n1337) );
  NAND4X1 U2287 ( .A(n1421), .B(n1422), .C(n1423), .D(n1424), .Q(
        n1419) );
  XNOR2X1 U2288 ( .A(g330), .B(g406), .Q(n1421) );
  XNOR2X1 U2289 ( .A(g309), .B(g416), .Q(n1422) );
  AO22X1 U2290 ( .A(g305), .B(n1910), .C(n1238), .D(n1903), .Q(n1221)
         );
  XNOR2X1 U2291 ( .A(n1240), .B(n1241), .Q(n1238) );
  NAND4X1 U2292 ( .A(n1884), .B(n1594), .C(n1646), .D(n1606), .Q(
        n1240) );
  AO221X1 U2293 ( .A(n1181), .B(g10720), .C(n1362), .D(g10724), .E(
        n1467), .Q(n1464) );
  AO222X1 U2294 ( .A(n1363), .B(n535), .C(g877), .D(n534), .E(n533), 
        .F(n532), .Q(n1467) );
  AO22X1 U2295 ( .A(g516), .B(n1902), .C(n1911), .D(g476), .Q(g11338)
         );
  AO22X1 U2296 ( .A(g506), .B(n1854), .C(g511), .D(n1911), .Q(g11336)
         );
  AO22X1 U2297 ( .A(g538), .B(n1854), .C(g534), .D(n1911), .Q(g11327)
         );
  AO22X1 U2298 ( .A(g530), .B(n1853), .C(g525), .D(n1913), .Q(g11329)
         );
  AO22X1 U2299 ( .A(g501), .B(n1902), .C(g506), .D(n1915), .Q(g11335)
         );
  AO22X1 U2300 ( .A(g525), .B(n1854), .C(g521), .D(n1913), .Q(g11330)
         );
  AO22X1 U2301 ( .A(n1241), .B(n1853), .C(g481), .D(n1914), .Q(g11324)
         );
  AO22X1 U2302 ( .A(g416), .B(n1902), .C(g421), .D(n1918), .Q(g11270)
         );
  AO22X1 U2303 ( .A(g486), .B(n1854), .C(g491), .D(n1912), .Q(g11332)
         );
  AO22X1 U2304 ( .A(g511), .B(n1853), .C(g516), .D(n1911), .Q(g11337)
         );
  AO22X1 U2305 ( .A(g496), .B(n1902), .C(g501), .D(n1912), .Q(g11334)
         );
  AO22X1 U2306 ( .A(g534), .B(n1853), .C(g530), .D(n1911), .Q(g11328)
         );
  AO22X1 U2307 ( .A(g476), .B(n1902), .C(g542), .D(n1915), .Q(g11325)
         );
  AO22X1 U2308 ( .A(g411), .B(n1854), .C(g416), .D(n1917), .Q(g11269)
         );
  AO22X1 U2309 ( .A(g542), .B(n1853), .C(g538), .D(n1916), .Q(g11326)
         );
  AO22X1 U2310 ( .A(g481), .B(n1902), .C(g486), .D(n1912), .Q(g11331)
         );
  AO22X1 U2311 ( .A(g391), .B(n1854), .C(g396), .D(n1918), .Q(g11265)
         );
  AO22X1 U2312 ( .A(g491), .B(n1853), .C(g496), .D(n1916), .Q(g11333)
         );
  AO22X1 U2313 ( .A(g440), .B(n1903), .C(g435), .D(n1920), .Q(g11261)
         );
  AO22X1 U2314 ( .A(g435), .B(n1903), .C(g431), .D(n1921), .Q(g11262)
         );
  AO22X1 U2315 ( .A(g406), .B(n1903), .C(g411), .D(n1917), .Q(g11268)
         );
  AO22X1 U2316 ( .A(g401), .B(n1903), .C(g406), .D(n1916), .Q(g11267)
         );
  AO22X1 U2317 ( .A(g386), .B(n1903), .C(g391), .D(n1918), .Q(g11264)
         );
  AO22X1 U2318 ( .A(g444), .B(n1903), .C(g440), .D(n1920), .Q(g11260)
         );
  AO22X1 U2319 ( .A(g452), .B(n1903), .C(g448), .D(n1910), .Q(g11258)
         );
  AO22X1 U2320 ( .A(g426), .B(n1903), .C(g386), .D(n1918), .Q(g11263)
         );
  AO22X1 U2321 ( .A(g396), .B(n1903), .C(g401), .D(n1919), .Q(g11266)
         );
  AO22X1 U2322 ( .A(g448), .B(n1903), .C(g444), .D(n1919), .Q(g11259)
         );
  AO22X1 U2323 ( .A(n602), .B(n1903), .C(g426), .D(n1914), .Q(g11256)
         );
  INVX1 U2324 ( .IN(n1390), .Q(n602) );
  AO22X1 U2325 ( .A(g421), .B(n1903), .C(g452), .D(n1921), .Q(g11257)
         );
  AO22X1 U2326 ( .A(g833), .B(n1855), .C(g947), .D(n1361), .Q(g11300)
         );
  AO22X1 U2327 ( .A(g845), .B(n1855), .C(g956), .D(n1361), .Q(g11306)
         );
  AO22X1 U2328 ( .A(g837), .B(n1855), .C(g950), .D(n1361), .Q(g11303)
         );
  AO22X1 U2329 ( .A(g861), .B(n1855), .C(g968), .D(n1361), .Q(g11314)
         );
  AO22X1 U2330 ( .A(g841), .B(n1855), .C(g953), .D(n1361), .Q(g11305)
         );
  AO22X1 U2331 ( .A(g829), .B(n1855), .C(g944), .D(n1361), .Q(g11298)
         );
  AO22X1 U2332 ( .A(g857), .B(n1855), .C(g965), .D(n1361), .Q(g11312)
         );
  AO22X1 U2333 ( .A(g853), .B(n1855), .C(g962), .D(n1361), .Q(g11310)
         );
  AO22X1 U2334 ( .A(g849), .B(n1855), .C(g959), .D(n1361), .Q(g11308)
         );
  AO22X1 U2335 ( .A(g339), .B(n1592), .C(n592), .D(n1244), .Q(g11478)
         );
  AO22X1 U2336 ( .A(g363), .B(n1592), .C(n592), .D(n1252), .Q(g11486)
         );
  AO22X1 U2337 ( .A(g351), .B(n1592), .C(n592), .D(n1247), .Q(g11482)
         );
  AO22X1 U2338 ( .A(g348), .B(n1592), .C(n592), .D(n1245), .Q(g11481)
         );
  AO22X1 U2339 ( .A(g366), .B(n1592), .C(n592), .D(n1253), .Q(g11487)
         );
  AO22X1 U2340 ( .A(g360), .B(n1592), .C(n592), .D(n1250), .Q(g11485)
         );
  AO22X1 U2341 ( .A(g342), .B(n1592), .C(n592), .D(n1254), .Q(g11488)
         );
  AO22X1 U2342 ( .A(g357), .B(n1592), .C(n592), .D(n1249), .Q(g11484)
         );
  AO22X1 U2343 ( .A(g354), .B(n1592), .C(n592), .D(n1248), .Q(g11483)
         );
  AO21X1 U2344 ( .A(g312), .B(n1907), .C(n1322), .Q(n1244) );
  OA221X1 U2345 ( .A(n1323), .B(g476), .C(n1599), .D(n1324), .E(
        n1854), .Q(n1322) );
  NAND2X1 U2346 ( .A(n610), .B(n674), .Q(n1324) );
  NOR2X1 U2347 ( .A(n1325), .B(n1306), .Q(n1323) );
  NOR2X1 U2348 ( .A(n1333), .B(n1334), .Q(g11393) );
  OA22X1 U2349 ( .A(n616), .B(n1335), .C(n1336), .D(n1722), .Q(n1333)
         );
  NOR2X1 U2350 ( .A(n1337), .B(n1338), .Q(n1336) );
  NOR2X1 U2351 ( .A(n1339), .B(n1334), .Q(g11392) );
  OA22X1 U2352 ( .A(n1340), .B(n1341), .C(n522), .D(n1720), .Q(n1339)
         );
  NAND2X1 U2353 ( .A(g976), .B(n1342), .Q(n1341) );
  NOR2X1 U2354 ( .A(n1343), .B(n1334), .Q(g11391) );
  XOR2X1 U2355 ( .A(n1340), .B(g976), .Q(n1343) );
  NOR2X1 U2356 ( .A(n1359), .B(n536), .Q(g11320) );
  XOR2X1 U2357 ( .A(g369), .B(n1360), .Q(n1359) );
  NOR2X1 U2358 ( .A(n1351), .B(n1334), .Q(g11349) );
  XOR2X1 U2359 ( .A(g971), .B(n1337), .Q(n1351) );
  OA21X1 U2360 ( .A(n1346), .B(n1347), .C(n521), .Q(g11376) );
  INVX1 U2361 ( .IN(n1345), .Q(n521) );
  OA21X1 U2362 ( .A(n1302), .B(n527), .C(g466), .Q(n1347) );
  NOR4X1 U2363 ( .A(n614), .B(n1594), .C(n1641), .D(n527), .Q(n1346)
         );
  OA21X1 U2364 ( .A(n1383), .B(g382), .C(n1384), .Q(g11292) );
  NOR2X1 U2365 ( .A(n1385), .B(n1360), .Q(n1383) );
  OA21X1 U2366 ( .A(n1386), .B(n1387), .C(n1384), .Q(g11291) );
  OA21X1 U2367 ( .A(n1385), .B(n1360), .C(g378), .Q(n1387) );
  AND4X1 U2368 ( .A(n1385), .B(g369), .C(g374), .D(n526), .Q(n1386) );
  NAND2X1 U2369 ( .A(n524), .B(g971), .Q(n1340) );
  NOR2X1 U2370 ( .A(n1388), .B(n536), .Q(g11290) );
  XOR2X1 U2371 ( .A(n1389), .B(g374), .Q(n1388) );
  AO22X1 U2372 ( .A(g1669), .B(n1888), .C(n1403), .D(n1404), .Q(g10865) );
  OA21X1 U2373 ( .A(g10722), .B(n1966), .C(n1875), .Q(n1403) );
  AO22X1 U2374 ( .A(n561), .B(n535), .C(g1730), .D(n1451), .Q(g10707)
         );
  AO22X1 U2375 ( .A(n1875), .B(n1452), .C(g1657), .D(n1888), .Q(g10767) );
  AO22X1 U2376 ( .A(g560), .B(n1930), .C(n1954), .D(n1405), .Q(g10797)
         );
  AO22X1 U2377 ( .A(g1681), .B(n1929), .C(n1955), .D(n1405), .Q(g10864) );
  AO22X1 U2378 ( .A(g572), .B(n1930), .C(n1954), .D(n1452), .Q(g10718)
         );
  AO221X1 U2379 ( .A(n1032), .B(n1364), .C(n619), .D(g1857), .E(
        n1365), .Q(g11294) );
  AND3X1 U2380 ( .A(n1366), .B(n1682), .C(n926), .Q(n1365) );
  NAND4X1 U2381 ( .A(n1367), .B(n1368), .C(n1369), .D(n1370), .Q(
        n1364) );
  NAND4X1 U2382 ( .A(n815), .B(n822), .C(n920), .D(n817), .Q(n1366)
         );
  AO22X1 U2383 ( .A(g1811), .B(n1054), .C(n555), .D(n1391), .Q(g10936)
         );
  NAND4X1 U2384 ( .A(n1291), .B(n547), .C(n535), .D(n1392), .Q(n1391)
         );
  AND3X1 U2385 ( .A(n545), .B(n544), .C(n546), .Q(n1392) );
  NAND4X1 U2386 ( .A(n1523), .B(n1524), .C(n1525), .D(n1526), .Q(
        g10720) );
  AOI222X1 U2387 ( .A(n1479), .B(g1552), .C(n572), .D(g1747), .E(
        n1480), .F(g1595), .Q(n1523) );
  AOI222X1 U2388 ( .A(n575), .B(g1724), .C(n578), .D(g4), .E(n579), 
        .F(g12), .Q(n1524) );
  OA221X1 U2389 ( .A(n583), .B(DFF_384_n1), .C(n577), .D(n1635), .E(
        n1532), .Q(n1525) );
  NOR3X1 U2390 ( .A(n1527), .B(n1528), .C(n1529), .Q(n1526) );
  AO222X1 U2391 ( .A(g953), .B(n580), .C(g932), .D(n1508), .E(g976), 
        .F(n1506), .Q(n1529) );
  NAND4X1 U2392 ( .A(n1558), .B(n1559), .C(n1560), .D(n1561), .Q(
        g10663) );
  NOR4X1 U2393 ( .A(n1562), .B(n1563), .C(n581), .D(n1564), .Q(n1561)
         );
  AOI22X1 U2394 ( .A(n572), .B(g1762), .C(n1483), .D(g281), .Q(n1558)
         );
  AOI222X1 U2395 ( .A(n1484), .B(n1637), .C(n1485), .D(g1586), .E(
        n1486), .F(g1543), .Q(n1560) );
  NAND4X1 U2396 ( .A(n1487), .B(n1488), .C(n1489), .D(n1490), .Q(
        g10724) );
  OA221X1 U2397 ( .A(n1494), .B(DFF_122_n1), .C(n1495), .D(DFF_445_n1), 
        .E(n1496), .Q(n1489) );
  AOI221X1 U2398 ( .A(n1483), .B(g275), .C(n1482), .D(g299), .E(
        n1497), .Q(n1488) );
  OA221X1 U2399 ( .A(n583), .B(DFF_350_n1), .C(n577), .D(n1636), .E(
        n1498), .Q(n1487) );
  NAND4X1 U2400 ( .A(n1514), .B(n1515), .C(n1516), .D(n1517), .Q(
        g10721) );
  OA22X1 U2401 ( .A(n577), .B(n1652), .C(n583), .D(DFF_242_n1), .Q(
        n1514) );
  AOI222X1 U2402 ( .A(n1485), .B(g1574), .C(n1482), .D(g293), .E(
        n1483), .F(g269), .Q(n1515) );
  AOI221X1 U2403 ( .A(n1479), .B(g1555), .C(n1480), .D(g1598), .E(
        n1522), .Q(n1516) );
  NAND4X1 U2404 ( .A(n1533), .B(n1534), .C(n1535), .D(n1536), .Q(
        g10719) );
  AOI222X1 U2405 ( .A(n1479), .B(g1549), .C(n572), .D(g1744), .E(
        n1480), .F(g1592), .Q(n1533) );
  OA221X1 U2406 ( .A(n583), .B(DFF_168_n1), .C(n577), .D(n1649), .E(
        n1549), .Q(n1535) );
  NAND4X1 U2407 ( .A(n1468), .B(n1469), .C(n1470), .D(n1471), .Q(
        g10726) );
  AOI222X1 U2408 ( .A(n1479), .B(g1564), .C(n572), .D(g1759), .E(
        n1480), .F(g1607), .Q(n1470) );
  AOI222X1 U2409 ( .A(n1484), .B(n1650), .C(n1485), .D(g1583), .E(
        n1486), .F(g1540), .Q(n1468) );
  OA221X1 U2410 ( .A(n1472), .B(n1638), .C(n1491), .D(n1492), .E(
        n1493), .Q(n1490) );
  NAND2X1 U2411 ( .A(n573), .B(n1477), .Q(n1492) );
  OA221X1 U2412 ( .A(n1472), .B(n1639), .C(n1473), .D(n1474), .E(
        n1475), .Q(n1471) );
  NAND2X1 U2413 ( .A(n1477), .B(n1478), .Q(n1474) );
  AO222X1 U2414 ( .A(n572), .B(g1750), .C(n579), .D(g9), .E(n575), 
        .F(g1727), .Q(n1522) );
  AO222X1 U2415 ( .A(g1333), .B(n576), .C(g1308), .D(n1511), .E(
        g4214), .F(n1476), .Q(n1562) );
  AO22X1 U2416 ( .A(n1480), .B(g1604), .C(n1479), .D(g1561), .Q(n1497)
         );
  AO22X1 U2417 ( .A(g4202), .B(n1481), .C(g944), .D(n1506), .Q(n1563)
         );
  ISOLANDX1 U2418 ( .D(g968), .ISO(n1472), .Q(n1564) );
  NOR4X1 U2419 ( .A(n1537), .B(n1538), .C(n1539), .D(n1540), .Q(n1536) );
  AO222X1 U2420 ( .A(g950), .B(n580), .C(g928), .D(n1508), .E(g971), 
        .F(n1506), .Q(n1539) );
  AO222X1 U2421 ( .A(g4204), .B(n1530), .C(g119), .D(n579), .E(g4191), .F(n1507), .Q(n1538) );
  NAND3X1 U2422 ( .A(n574), .B(n1541), .C(n1542), .Q(n1537) );
  NAND2X1 U2423 ( .A(g123), .B(n578), .Q(n1542) );
  INVX1 U2424 ( .IN(n1509), .Q(n574) );
  NOR3X1 U2425 ( .A(n1518), .B(n1519), .C(n1520), .Q(n1517) );
  AO222X1 U2426 ( .A(g981), .B(n1506), .C(g956), .D(n580), .E(g4198), 
        .F(n1481), .Q(n1520) );
  AOI22X1 U2427 ( .A(g4200), .B(n1481), .C(g1580), .D(n1485), .Q(
        n1498) );
  AOI22X1 U2428 ( .A(n575), .B(g1733), .C(n572), .D(g1756), .Q(n1496)
         );
  AOI222X1 U2429 ( .A(n1485), .B(g1567), .C(n1482), .D(g287), .E(
        n1483), .F(g263), .Q(n1549) );
  OA22X1 U2430 ( .A(n1543), .B(n1568), .C(n1550), .D(n1640), .Q(n1559)
         );
  NAND2X1 U2431 ( .A(n573), .B(n1478), .Q(n1568) );
  NAND2X1 U2432 ( .A(g1317), .B(n550), .Q(n1255) );
  NAND3X1 U2433 ( .A(n1113), .B(n1270), .C(n629), .Q(n1227) );
  NAND4X1 U2434 ( .A(n1271), .B(n1272), .C(n1273), .D(n1274), .Q(
        n1270) );
  XNOR2X1 U2435 ( .A(test_so2), .B(g1255), .Q(n1271) );
  XNOR2X1 U2436 ( .A(g1015), .B(g1265), .Q(n1272) );
  AO21X1 U2437 ( .A(g201), .B(n1880), .C(n1288), .Q(n1261) );
  OA221X1 U2438 ( .A(n1289), .B(n1699), .C(n627), .D(n1290), .E(
        n1959), .Q(n1288) );
  INVX1 U2439 ( .IN(n1289), .Q(n627) );
  AO22X1 U2440 ( .A(g1766), .B(n1653), .C(n1882), .D(g10719), .Q(n1373) );
  AO22X1 U2441 ( .A(g1776), .B(n1653), .C(n1882), .D(g10721), .Q(n1374) );
  AO22X1 U2442 ( .A(n1862), .B(n1863), .C(n1864), .D(g1280), .Q(n1326)
         );
  OAI21X1 U2443 ( .A(n1328), .B(n1329), .C(n1864), .Q(n1863) );
  INVX1 U2444 ( .IN(g109), .Q(n1988) );
  INVX1 U2445 ( .IN(g109), .Q(n1987) );
  AO22X1 U2446 ( .A(n549), .B(g1791), .C(g1324), .D(n1255), .Q(g11607)
         );
  AO22X1 U2447 ( .A(n549), .B(g1776), .C(g1314), .D(n1255), .Q(g11604)
         );
  AO22X1 U2448 ( .A(n549), .B(g1781), .C(g1318), .D(n1255), .Q(g11605)
         );
  AO22X1 U2449 ( .A(n549), .B(g1796), .C(g1327), .D(n1255), .Q(g11608)
         );
  AO22X1 U2450 ( .A(n549), .B(g1786), .C(g1321), .D(n1255), .Q(g11606)
         );
  AO22X1 U2451 ( .A(g546), .B(n1925), .C(n1954), .D(n1412), .Q(g10791)
         );
  AO22X1 U2452 ( .A(g575), .B(n1927), .C(n1954), .D(n1411), .Q(g10800)
         );
  AO22X1 U2453 ( .A(g557), .B(n1926), .C(n1954), .D(n1408), .Q(g10795)
         );
  AO22X1 U2454 ( .A(g549), .B(n1927), .C(n1954), .D(n1409), .Q(g10855)
         );
  AO22X1 U2455 ( .A(g1678), .B(n1929), .C(n1955), .D(n1408), .Q(g10862) );
  AO22X1 U2456 ( .A(g1675), .B(n1928), .C(n1955), .D(n1410), .Q(g10860) );
  AO22X1 U2457 ( .A(g554), .B(n1926), .C(n1954), .D(n1410), .Q(g10793)
         );
  AO22X1 U2458 ( .A(g1672), .B(n1928), .C(n1954), .D(n1412), .Q(g10858) );
  AO22X1 U2459 ( .A(g1666), .B(n1888), .C(n1406), .D(n1875), .Q(g10863) );
  OA21X1 U2460 ( .A(n532), .B(g1718), .C(n1407), .Q(n1406) );
  AO22X1 U2461 ( .A(n549), .B(test_so5), .C(test_so9), .D(n1255), .Q(
        g11603) );
  AO22X1 U2462 ( .A(n549), .B(g1801), .C(g1330), .D(n1255), .Q(g11609)
         );
  AO22X1 U2463 ( .A(n549), .B(g1806), .C(g1333), .D(n1255), .Q(g11610)
         );
  AO22X1 U2464 ( .A(n549), .B(g1766), .C(g1308), .D(n1255), .Q(g11602)
         );
  AO22X1 U2465 ( .A(g1663), .B(n1888), .C(n1875), .D(n1409), .Q(g10861) );
  AO22X1 U2466 ( .A(g1660), .B(n1888), .C(n1875), .D(n1411), .Q(g10859) );
  AO221X1 U2467 ( .A(test_so5), .B(n1373), .C(g1781), .D(n1374), .E(
        n1881), .Q(n1368) );
  ISOLANDX1 U2468 ( .D(g1336), .ISO(n1227), .Q(n1231) );
  NOR2X1 U2469 ( .A(n1223), .B(n1224), .Q(g11641) );
  OA22X1 U2470 ( .A(n687), .B(n1225), .C(n1226), .D(n1721), .Q(n1223)
         );
  NOR2X1 U2471 ( .A(n1227), .B(n1228), .Q(n1226) );
  NOR2X1 U2472 ( .A(n1233), .B(n1224), .Q(g11639) );
  XNOR2X1 U2473 ( .A(g1341), .B(n1231), .Q(n1233) );
  NOR2X1 U2474 ( .A(n1234), .B(n1224), .Q(g11636) );
  XOR2X1 U2475 ( .A(n1227), .B(g1336), .Q(n1234) );
  NOR2X1 U2476 ( .A(n1230), .B(n1224), .Q(g11640) );
  AOI22X1 U2477 ( .A(n1231), .B(n1232), .C(n1225), .D(g1346), .Q(
        n1230) );
  ISOLANDX1 U2478 ( .D(g1341), .ISO(n1229), .Q(n1232) );
  XNOR2X1 U2479 ( .A(n1332), .B(g1027), .Q(n1285) );
  NAND2X1 U2480 ( .A(g1032), .B(n1222), .Q(n1332) );
  NOR3X1 U2481 ( .A(n1281), .B(n1282), .C(n1283), .Q(n1273) );
  XOR2X1 U2482 ( .A(test_so6), .B(g1023), .Q(n1281) );
  XOR2X1 U2483 ( .A(g1260), .B(g1019), .Q(n1283) );
  XOR2X1 U2484 ( .A(n1284), .B(n1285), .Q(n1282) );
  AO22X1 U2485 ( .A(g1618), .B(n1930), .C(n1955), .D(n1256), .Q(g11579) );
  XOR2X1 U2486 ( .A(g1610), .B(n1257), .Q(n1256) );
  OA22X1 U2487 ( .A(n1258), .B(n1259), .C(n1260), .D(n1261), .Q(n1257)
         );
  ISOLANDX1 U2488 ( .D(n1262), .ISO(n1258), .Q(n1260) );
  OAI22X1 U2489 ( .A(n1375), .B(n715), .C(n1032), .D(n1376), .Q(
        g11293) );
  OA21X1 U2490 ( .A(n1377), .B(DFF_311_n1), .C(n815), .Q(n1376) );
  OA22X1 U2491 ( .A(g10719), .B(n1653), .C(g1806), .D(n1882), .Q(n1375) );
  AND3X1 U2492 ( .A(n1378), .B(n1379), .C(g4904), .Q(n1377) );
  AND3X1 U2493 ( .A(n1956), .B(n1610), .C(g1289), .Q(n1113) );
  INVX1 U2494 ( .IN(n1924), .Q(n1956) );
  NOR3X1 U2495 ( .A(n1983), .B(n1865), .C(n1866), .Q(n1362) );
  NAND3X1 U2496 ( .A(n1977), .B(DFF_121_n1), .C(g2986), .Q(n1059) );
  NAND3X1 U2497 ( .A(n1977), .B(DFF_194_n1), .C(g3069), .Q(n1236) );
  AO22X1 U2498 ( .A(g1796), .B(n1653), .C(n1882), .D(g10663), .Q(n1372) );
  AO22X1 U2499 ( .A(g1786), .B(n1653), .C(n1882), .D(g10724), .Q(n1371) );
  OR2X1 U2500 ( .A(n1484), .B(g6254), .Q(n1867) );
  AO22X1 U2501 ( .A(g1275), .B(n1113), .C(g1235), .D(n1120), .Q(g7296)
         );
  AO22X1 U2502 ( .A(g1304), .B(n1113), .C(g1300), .D(n1120), .Q(g7291)
         );
  AO22X1 U2503 ( .A(g1292), .B(n1113), .C(g1284), .D(n1120), .Q(g7294)
         );
  AO22X1 U2504 ( .A(g1255), .B(n1113), .C(g1260), .D(n1120), .Q(g7301)
         );
  AO22X1 U2505 ( .A(g1284), .B(n1113), .C(g1280), .D(n1120), .Q(g7295)
         );
  AO22X1 U2506 ( .A(g1250), .B(n1113), .C(g1255), .D(n1120), .Q(g7300)
         );
  AO22X1 U2507 ( .A(g1240), .B(n1113), .C(g1245), .D(n1120), .Q(g7298)
         );
  AO22X1 U2508 ( .A(g1265), .B(n1113), .C(test_so6), .D(n1120), .Q(
        g7303) );
  AO22X1 U2509 ( .A(g1296), .B(n1113), .C(g1292), .D(n1120), .Q(g7293)
         );
  AO22X1 U2510 ( .A(g1245), .B(n1113), .C(g1250), .D(n1120), .Q(g7299)
         );
  AO22X1 U2511 ( .A(g1235), .B(n1113), .C(g1240), .D(n1120), .Q(g7297)
         );
  AO22X1 U2512 ( .A(g1300), .B(n1113), .C(g1296), .D(n1120), .Q(g7292)
         );
  AO22X1 U2513 ( .A(g1260), .B(n1113), .C(g1265), .D(n1120), .Q(g7302)
         );
  AO22X1 U2514 ( .A(test_so6), .B(n1113), .C(g1304), .D(n1120), .Q(
        g7290) );
  AO22X1 U2515 ( .A(g105), .B(n1930), .C(n1955), .D(n1393), .Q(g10898)
         );
  NAND2X1 U2516 ( .A(n1394), .B(n1222), .Q(n1393) );
  XOR3X1 U2517 ( .A(n1397), .B(n1398), .C(n1399), .Q(n1394) );
  XNOR2X1 U2518 ( .A(g1023), .B(g1027), .Q(n1399) );
  AO22X1 U2519 ( .A(n1875), .B(n1453), .C(g1654), .D(n1888), .Q(g10765) );
  AO22X1 U2520 ( .A(g1724), .B(n1451), .C(n528), .D(n561), .Q(g10771)
         );
  INVX1 U2521 ( .IN(n1414), .Q(n528) );
  AO22X1 U2522 ( .A(n1113), .B(n1284), .C(g1275), .D(n1120), .Q(g11443) );
  AO22X1 U2523 ( .A(g569), .B(n1928), .C(n1955), .D(n1453), .Q(g10717)
         );
  AO22X1 U2524 ( .A(g1687), .B(n1925), .C(n1954), .D(n1417), .Q(g10776) );
  AO22X1 U2525 ( .A(g566), .B(n1927), .C(n1954), .D(n1417), .Q(g10799)
         );
  AO22X1 U2526 ( .A(g563), .B(n1927), .C(n1954), .D(n1402), .Q(g10798)
         );
  AO22X1 U2527 ( .A(g1684), .B(n1929), .C(n1955), .D(n1402), .Q(g10866) );
  AO22X1 U2528 ( .A(g1733), .B(n1451), .C(n561), .D(n1382), .Q(g10711)
         );
  AO22X1 U2529 ( .A(n561), .B(n532), .C(g1727), .D(n1451), .Q(g10773)
         );
  AO22X1 U2530 ( .A(n561), .B(n534), .C(g1721), .D(n1451), .Q(g10770)
         );
  AO221X1 U2531 ( .A(g1791), .B(n1371), .C(g1801), .D(n1372), .E(
        n1882), .Q(n1370) );
  NOR2X1 U2532 ( .A(n1868), .B(n1967), .Q(n1363) );
  ISOLANDX1 U2533 ( .D(g178), .ISO(n1966), .Q(g6786) );
  ISOLANDX1 U2534 ( .D(g1424), .ISO(n1967), .Q(g6234) );
  AO21X1 U2535 ( .A(g123), .B(n1968), .C(n1132), .Q(g7032) );
  NOR4X1 U2536 ( .A(n1133), .B(n1134), .C(n1135), .D(n1136), .Q(n1132) );
  OR4X1 U2537 ( .A(g148), .B(g153), .C(g158), .D(g162), .Q(n1133) );
  OR4X1 U2538 ( .A(g131), .B(g135), .C(g139), .D(g143), .Q(n1134) );
  INVX1 U2539 ( .IN(g1703), .Q(n744) );
  OA21X1 U2540 ( .A(n1107), .B(n1108), .C(n1109), .Q(g7586) );
  OA21X1 U2541 ( .A(n1110), .B(n1103), .C(g1227), .Q(n1108) );
  AND4X1 U2542 ( .A(n1110), .B(g1218), .C(g1223), .D(n557), .Q(n1107)
         );
  NOR2X1 U2543 ( .A(n1965), .B(n1286), .Q(g11514) );
  XOR3X1 U2544 ( .A(n1261), .B(g1415), .C(n1287), .Q(n1286) );
  XOR3X1 U2545 ( .A(g1515), .B(g1448), .C(n1602), .Q(n1287) );
  AO22X1 U2546 ( .A(g1), .B(n1975), .C(n1154), .D(n1155), .Q(g6679) );
  NOR2X1 U2547 ( .A(n1156), .B(n1157), .Q(n1155) );
  NOR4X1 U2548 ( .A(n1158), .B(n1710), .C(n1602), .D(n1627), .Q(n1154) );
  OR4X1 U2549 ( .A(g1403), .B(g1407), .C(g1411), .D(g1415), .Q(n1156)
         );
  XNOR2X1 U2550 ( .A(n1381), .B(n1382), .Q(n1378) );
  OA22X1 U2551 ( .A(g1857), .B(n1380), .C(n1682), .D(n920), .Q(n1381)
         );
  OR2X1 U2552 ( .A(g845), .B(g849), .Q(n1443) );
  NAND4X1 U2553 ( .A(g6234), .B(n1159), .C(g1432), .D(g1448), .Q(
        n1158) );
  NOR2X1 U2554 ( .A(n1111), .B(n540), .Q(g7581) );
  XOR2X1 U2555 ( .A(n1112), .B(g1223), .Q(n1111) );
  NAND2X1 U2556 ( .A(n557), .B(g1218), .Q(n1112) );
  NOR2X1 U2557 ( .A(n1102), .B(n540), .Q(g7632) );
  XOR2X1 U2558 ( .A(n1103), .B(g1218), .Q(n1102) );
  NAND4X1 U2559 ( .A(g182), .B(g6786), .C(n1137), .D(g166), .Q(n1136)
         );
  NOR2X1 U2560 ( .A(n1106), .B(n540), .Q(g7590) );
  AOI21X1 U2561 ( .A(n665), .B(n557), .C(g1231), .Q(n1106) );
  INVX1 U2562 ( .IN(n1724), .Q(n560) );
  AO22X1 U2563 ( .A(g1687), .B(n1882), .C(g1669), .D(n1653), .Q(g6955)
         );
  AO22X1 U2564 ( .A(g1684), .B(n1882), .C(g1666), .D(n1653), .Q(g6949)
         );
  AO22X1 U2565 ( .A(g1681), .B(n1882), .C(g1663), .D(n1653), .Q(g6942)
         );
  AO22X1 U2566 ( .A(g1678), .B(n1882), .C(g1660), .D(n1653), .Q(g6932)
         );
  AO22X1 U2567 ( .A(g1675), .B(n1882), .C(g1657), .D(n1653), .Q(g6926)
         );
  AO22X1 U2568 ( .A(g1672), .B(n1882), .C(g1654), .D(n1653), .Q(g6920)
         );
  AO21X1 U2569 ( .A(g617), .B(n959), .C(n960), .Q(n899) );
  AO21X1 U2570 ( .A(g1840), .B(n926), .C(n929), .Q(n853) );
  NAND4X1 U2571 ( .A(n1184), .B(n1185), .C(n1186), .D(n1187), .Q(
        n1183) );
  NOR4X1 U2572 ( .A(n1188), .B(g192), .C(g248), .D(g197), .Q(n1187)
         );
  AND3X1 U2573 ( .A(n1977), .B(n1700), .C(g201), .Q(n1186) );
  NAND3X1 U2574 ( .A(n1711), .B(n1629), .C(n1603), .Q(n1188) );
  NAND2X1 U2575 ( .A(g1765), .B(g1610), .Q(n1217) );
  NAND2X1 U2576 ( .A(n1137), .B(n1613), .Q(n1145) );
  NOR2X1 U2577 ( .A(n1964), .B(test_so1), .Q(n1046) );
  NOR2X1 U2578 ( .A(n1724), .B(g4089), .Q(g6842) );
  AO22X1 U2579 ( .A(g673), .B(n899), .C(n648), .D(n914), .Q(n913) );
  XOR2X1 U2580 ( .A(g658), .B(n718), .Q(n914) );
  AO22X1 U2581 ( .A(g1887), .B(n853), .C(n622), .D(n871), .Q(n870) );
  XOR2X1 U2582 ( .A(g1872), .B(n712), .Q(n871) );
  NOR2X1 U2583 ( .A(n892), .B(g1891), .Q(n877) );
  NOR2X1 U2584 ( .A(n950), .B(g677), .Q(n935) );
  NAND2X1 U2585 ( .A(g1104), .B(n985), .Q(n978) );
  NAND2X1 U2586 ( .A(g461), .B(n1641), .Q(n1306) );
  NOR2X1 U2587 ( .A(n662), .B(g1718), .Q(n1404) );
  OA21X1 U2588 ( .A(n1609), .B(g591), .C(n668), .Q(n1160) );
  OA21X1 U2589 ( .A(n1655), .B(g1814), .C(n715), .Q(n1148) );
  NAND2X1 U2590 ( .A(g599), .B(n1593), .Q(n953) );
  NAND2X1 U2591 ( .A(g599), .B(n1607), .Q(n1025) );
  NAND2X1 U2592 ( .A(g1822), .B(n1608), .Q(n920) );
  AO21X1 U2593 ( .A(g869), .B(n1352), .C(n1966), .Q(n1334) );
  NAND2X1 U2594 ( .A(n1724), .B(n744), .Q(n1054) );
  NAND2X1 U2595 ( .A(n1970), .B(DFF_441_n1), .Q(n1345) );
  NOR2X1 U2596 ( .A(n1965), .B(g869), .Q(n1384) );
  AND3X1 U2597 ( .A(g743), .B(n1969), .C(g744), .Q(g5659) );
  AND3X1 U2598 ( .A(g741), .B(n1976), .C(g742), .Q(g5658) );
  NAND2X1 U2599 ( .A(g4180), .B(n1093), .Q(n1092) );
  NAND2X1 U2600 ( .A(g466), .B(n1606), .Q(n1307) );
  NOR3X1 U2601 ( .A(g591), .B(g611), .C(n964), .Q(n954) );
  NAND2X1 U2602 ( .A(g471), .B(n1646), .Q(n1325) );
  NOR2X1 U2603 ( .A(n1962), .B(g1212), .Q(n1109) );
  NAND2X1 U2604 ( .A(g591), .B(n1644), .Q(n966) );
  NAND2X1 U2605 ( .A(g627), .B(n1612), .Q(n1119) );
  NOR2X1 U2606 ( .A(n1966), .B(g1718), .Q(n1416) );
  NOR4X1 U2607 ( .A(n1654), .B(g1104), .C(g1107), .D(g1110), .Q(n1263) );
  NOR2X1 U2608 ( .A(n1614), .B(g1110), .Q(n985) );
  NAND3X1 U2609 ( .A(g745), .B(n1976), .C(g746), .Q(n1042) );
  NOR3X1 U2610 ( .A(g1814), .B(g1834), .C(n928), .Q(n1032) );
  NAND2X1 U2611 ( .A(g1231), .B(n665), .Q(n1114) );
  NAND3X1 U2612 ( .A(n1884), .B(g461), .C(g466), .Q(n1302) );
  NAND3X1 U2613 ( .A(n1614), .B(n1677), .C(g1104), .Q(n993) );
  NAND3X1 U2614 ( .A(n1646), .B(n1606), .C(g461), .Q(n1318) );
  NAND3X1 U2615 ( .A(test_so5), .B(g1766), .C(g1776), .Q(n1172) );
  NAND3X1 U2616 ( .A(n1658), .B(n1614), .C(g1110), .Q(n999) );
  NAND2X1 U2617 ( .A(g219), .B(g2355), .Q(n974) );
  NAND2X1 U2618 ( .A(g231), .B(g2355), .Q(n995) );
  NAND2X1 U2619 ( .A(g207), .B(g2355), .Q(n1001) );
  NAND2X1 U2620 ( .A(g225), .B(n1880), .Q(n981) );
  NAND2X1 U2621 ( .A(g186), .B(n1880), .Q(n989) );
  NAND2X1 U2622 ( .A(g237), .B(n1880), .Q(n1007) );
  NAND2X1 U2623 ( .A(g213), .B(n1880), .Q(n1012) );
  NAND2X1 U2624 ( .A(g1504), .B(n1969), .Q(n1166) );
  NAND2X1 U2625 ( .A(n1969), .B(DFF_126_n1), .Q(n1216) );
  NAND2X1 U2626 ( .A(g4174), .B(g4173), .Q(n1214) );
  NOR3X1 U2627 ( .A(g650), .B(g654), .C(n1128), .Q(n959) );
  NAND2X1 U2628 ( .A(g1828), .B(g1814), .Q(n817) );
  AND4X1 U2629 ( .A(n1845), .B(n1843), .C(n1847), .D(n799), .Q(n795)
         );
  NOR2X1 U2630 ( .A(g6258), .B(g6257), .Q(n799) );
  AO21X1 U2631 ( .A(n605), .B(n930), .C(n606), .Q(g8920) );
  XNOR2X1 U2632 ( .A(g713), .B(n931), .Q(n930) );
  NAND2X1 U2633 ( .A(n850), .B(n932), .Q(n931) );
  AO222X1 U2634 ( .A(n933), .B(n934), .C(n935), .D(n936), .E(g718), 
        .F(n899), .Q(n932) );
  NAND2X1 U2635 ( .A(g1814), .B(n1643), .Q(n826) );
  NAND2X1 U2636 ( .A(g1822), .B(n1605), .Q(n822) );
  NAND2X1 U2637 ( .A(g668), .B(n913), .Q(n912) );
  NAND2X1 U2638 ( .A(g1882), .B(n870), .Q(n869) );
  ISOLANDX1 U2639 ( .D(n962), .ISO(n958), .Q(n804) );
  OAI22X1 U2640 ( .A(n1696), .B(n902), .C(n901), .D(g731), .Q(n962)
         );
  ISOLANDX1 U2641 ( .D(n1147), .ISO(g1868), .Q(n926) );
  NAND3X1 U2642 ( .A(g1223), .B(g1218), .C(g1227), .Q(n1110) );
  NAND3X1 U2643 ( .A(n1607), .B(n1644), .C(g605), .Q(n832) );
  AND4X1 U2644 ( .A(n1624), .B(n1687), .C(n1206), .D(n1207), .Q(n1185)
         );
  NOR2X1 U2645 ( .A(g1386), .B(g1383), .Q(n1206) );
  NOR4X1 U2646 ( .A(g219), .B(g213), .C(g207), .D(g186), .Q(n1207) );
  NAND2X1 U2647 ( .A(g4176), .B(n1193), .Q(n1153) );
  NAND2X1 U2648 ( .A(g4178), .B(n1125), .Q(n1099) );
  AND4X1 U2649 ( .A(n936), .B(n1615), .C(n965), .D(n1662), .Q(n907) );
  NOR2X1 U2650 ( .A(g713), .B(g677), .Q(n965) );
  AND4X1 U2651 ( .A(n878), .B(n1616), .C(n919), .D(n1663), .Q(n862) );
  NOR2X1 U2652 ( .A(g1927), .B(g1891), .Q(n919) );
  NAND2X1 U2653 ( .A(g798), .B(g794), .Q(n1029) );
  ISOLANDX1 U2654 ( .D(g746), .ISO(g750), .Q(g4171) );
  NAND3X1 U2655 ( .A(n959), .B(n1609), .C(g617), .Q(n1016) );
  NAND3X1 U2656 ( .A(n926), .B(n1655), .C(g1840), .Q(n1031) );
  NOR2X1 U2657 ( .A(g611), .B(n834), .Q(n1024) );
  ISOLANDX1 U2658 ( .D(n917), .ISO(n918), .Q(n812) );
  OAI22X1 U2659 ( .A(n1697), .B(n857), .C(n856), .D(g1945), .Q(n917)
         );
  AND3X1 U2660 ( .A(g1909), .B(g1900), .C(g1918), .Q(n876) );
  AND3X1 U2661 ( .A(g695), .B(g686), .C(g704), .Q(n934) );
  NAND2X1 U2662 ( .A(n1007), .B(n1008), .Q(n969) );
  AO221X1 U2663 ( .A(n1009), .B(g1145), .C(n1617), .D(n1010), .E(
        g2355), .Q(n1008) );
  NOR2X1 U2664 ( .A(n999), .B(n1654), .Q(n1009) );
  NAND2X1 U2665 ( .A(g1101), .B(n634), .Q(n1010) );
  NAND2X1 U2666 ( .A(n1012), .B(n1013), .Q(n979) );
  AO221X1 U2667 ( .A(n1014), .B(g1129), .C(n1705), .D(n1015), .E(
        n1880), .Q(n1013) );
  NAND2X1 U2668 ( .A(n633), .B(g1101), .Q(n1015) );
  NOR2X1 U2669 ( .A(n1654), .B(n1005), .Q(n1014) );
  NAND2X1 U2670 ( .A(n1001), .B(n1002), .Q(n986) );
  AO221X1 U2671 ( .A(n1003), .B(g1125), .C(n1708), .D(n1004), .E(
        n1880), .Q(n1002) );
  NAND2X1 U2672 ( .A(n633), .B(n1654), .Q(n1004) );
  NOR2X1 U2673 ( .A(g1101), .B(n1005), .Q(n1003) );
  NAND2X1 U2674 ( .A(n974), .B(n975), .Q(n973) );
  AO221X1 U2675 ( .A(n976), .B(g1133), .C(n1706), .D(n977), .E(n1880), .Q(n975) );
  NAND2X1 U2676 ( .A(n631), .B(n1654), .Q(n977) );
  NOR2X1 U2677 ( .A(g1101), .B(n978), .Q(n976) );
  NOR2X1 U2678 ( .A(g4173), .B(n537), .Q(g4940) );
  NAND2X1 U2679 ( .A(g4181), .B(n630), .Q(n1045) );
  AO22X1 U2680 ( .A(g192), .B(n1880), .C(g1512), .D(n1959), .Q(n1082)
         );
  AO22X1 U2681 ( .A(g243), .B(n1880), .C(g1633), .D(n1959), .Q(n1069)
         );
  AO22X1 U2682 ( .A(g248), .B(g2355), .C(g1636), .D(n1959), .Q(n1077)
         );
  ISOLANDX1 U2683 ( .D(g382), .ISO(n1385), .Q(n1420) );
  AO22X1 U2684 ( .A(g192), .B(g2355), .C(g549), .D(n1959), .Q(g6049)
         );
  AO22X1 U2685 ( .A(g248), .B(n1880), .C(g575), .D(n1959), .Q(g6045)
         );
  AO22X1 U2686 ( .A(g243), .B(g2355), .C(g572), .D(n1959), .Q(g6042)
         );
  AO21X1 U2687 ( .A(n805), .B(n963), .C(n649), .Q(n958) );
  NAND2X1 U2688 ( .A(g639), .B(n964), .Q(n963) );
  NAND4X1 U2689 ( .A(n648), .B(g668), .C(g658), .D(n908), .Q(n949) );
  NAND4X1 U2690 ( .A(n622), .B(g1882), .C(g1872), .D(n863), .Q(n891)
         );
  AO21X1 U2691 ( .A(g1639), .B(n1922), .C(n1049), .Q(g8193) );
  OA221X1 U2692 ( .A(n1050), .B(test_so4), .C(n1661), .D(n1051), .E(
        n1953), .Q(n1049) );
  NAND2X1 U2693 ( .A(n632), .B(n1654), .Q(n1051) );
  NOR2X1 U2694 ( .A(g1101), .B(n993), .Q(n1050) );
  AND3X1 U2695 ( .A(n831), .B(n832), .C(n833), .Q(n829) );
  NAND2X1 U2696 ( .A(n834), .B(g599), .Q(n833) );
  OA221X1 U2697 ( .A(n806), .B(g1834), .C(n623), .D(n807), .E(g2355), 
        .Q(g9555) );
  NAND2X1 U2698 ( .A(g1834), .B(n808), .Q(n807) );
  ISOLANDX1 U2699 ( .D(n808), .ISO(n623), .Q(n806) );
  AO21X1 U2700 ( .A(n809), .B(n598), .C(g1840), .Q(n808) );
  AND3X1 U2701 ( .A(n1044), .B(n1045), .C(n1046), .Q(g8244) );
  OR2X1 U2702 ( .A(g4181), .B(n630), .Q(n1044) );
  AND3X1 U2703 ( .A(n1215), .B(n1214), .C(n1046), .Q(g5529) );
  OR2X1 U2704 ( .A(g4173), .B(g4174), .Q(n1215) );
  AND3X1 U2705 ( .A(n1192), .B(n1153), .C(n1046), .Q(g6123) );
  OR2X1 U2706 ( .A(g4176), .B(n1193), .Q(n1192) );
  AND3X1 U2707 ( .A(n1124), .B(n1099), .C(n1046), .Q(g7191) );
  OR2X1 U2708 ( .A(g4178), .B(n1125), .Q(n1124) );
  AND3X1 U2709 ( .A(n1091), .B(n1092), .C(n1046), .Q(g8019) );
  OR2X1 U2710 ( .A(n1093), .B(g4180), .Q(n1091) );
  AND3X1 U2711 ( .A(n1122), .B(n1097), .C(n520), .Q(g7202) );
  OR2X1 U2712 ( .A(g814), .B(n1123), .Q(n1122) );
  AND3X1 U2713 ( .A(n1190), .B(n1151), .C(n520), .Q(g6126) );
  OR2X1 U2714 ( .A(g806), .B(n1191), .Q(n1190) );
  AND3X1 U2715 ( .A(n1089), .B(n1043), .C(n520), .Q(g8024) );
  OR2X1 U2716 ( .A(n1090), .B(g822), .Q(n1089) );
  AND3X1 U2717 ( .A(n1149), .B(n1634), .C(n1977), .Q(g6747) );
  NAND2X1 U2718 ( .A(n1714), .B(DFF_452_n1), .Q(n1149) );
  NOR4X1 U2719 ( .A(n1203), .B(n1204), .C(g192), .D(g1400), .Q(n1202)
         );
  NAND3X1 U2720 ( .A(n1619), .B(n1598), .C(n1678), .Q(n1204) );
  NAND4X1 U2721 ( .A(n1184), .B(n1185), .C(n1205), .D(n1700), .Q(
        n1203) );
  NOR2X1 U2722 ( .A(g1397), .B(g1389), .Q(n1205) );
  NAND3X1 U2723 ( .A(g1786), .B(n1141), .C(g1791), .Q(n1117) );
  OAI22X1 U2724 ( .A(g1153), .B(n1685), .C(g1149), .D(n1265), .Q(
        n1264) );
  OA21X1 U2725 ( .A(n1266), .B(n1267), .C(n1686), .Q(n1265) );
  NAND4X1 U2726 ( .A(n1660), .B(n1617), .C(n1597), .D(n1269), .Q(
        n1266) );
  NAND4X1 U2727 ( .A(n1661), .B(n1618), .C(n1596), .D(n1268), .Q(
        n1267) );
  OR4X1 U2728 ( .A(n826), .B(g1828), .C(g1834), .D(g1840), .Q(n1038)
         );
  NAND2X1 U2729 ( .A(n926), .B(n927), .Q(n918) );
  AO21X1 U2730 ( .A(g1857), .B(n928), .C(n809), .Q(n927) );
  NAND3X1 U2731 ( .A(n1608), .B(n1643), .C(g1828), .Q(n815) );
  AO21X1 U2732 ( .A(g1627), .B(n1959), .C(n568), .Q(n1086) );
  AO21X1 U2733 ( .A(g1630), .B(n1958), .C(n569), .Q(n1088) );
  AO22X1 U2734 ( .A(g1415), .B(n1169), .C(n538), .D(g1567), .Q(g6468)
         );
  AO22X1 U2735 ( .A(g1466), .B(n1167), .C(n539), .D(g1555), .Q(g6534)
         );
  AO22X1 U2736 ( .A(g1504), .B(n1167), .C(n539), .D(g1528), .Q(g6522)
         );
  AO22X1 U2737 ( .A(g1448), .B(n1169), .C(n538), .D(g1607), .Q(g6515)
         );
  AO22X1 U2738 ( .A(g1407), .B(n1169), .C(n538), .D(g1586), .Q(g6514)
         );
  AO22X1 U2739 ( .A(g1470), .B(n1167), .C(n539), .D(g1552), .Q(g6529)
         );
  AO22X1 U2740 ( .A(g1436), .B(n1169), .C(n538), .D(g1598), .Q(g6481)
         );
  AO22X1 U2741 ( .A(g1474), .B(n1167), .C(n539), .D(g1549), .Q(g6523)
         );
  AO22X1 U2742 ( .A(g1490), .B(n1167), .C(n539), .D(g1537), .Q(g6537)
         );
  AO22X1 U2743 ( .A(g1432), .B(n1169), .C(n538), .D(g1595), .Q(g6479)
         );
  AO22X1 U2744 ( .A(g1419), .B(n1169), .C(n538), .D(g1577), .Q(g6480)
         );
  AO22X1 U2745 ( .A(g1508), .B(n1167), .C(n539), .D(g1524), .Q(g6513)
         );
  AO22X1 U2746 ( .A(g1403), .B(n1169), .C(n538), .D(g1592), .Q(g6470)
         );
  AO22X1 U2747 ( .A(g1486), .B(n1167), .C(n539), .D(g1540), .Q(g6541)
         );
  AO22X1 U2748 ( .A(g1478), .B(n1167), .C(n539), .D(g1546), .Q(g6551)
         );
  AO22X1 U2749 ( .A(g1458), .B(n1167), .C(n539), .D(g1561), .Q(g6542)
         );
  AO22X1 U2750 ( .A(g1424), .B(n1169), .C(n538), .D(g1583), .Q(g6506)
         );
  AO22X1 U2751 ( .A(g1440), .B(n1169), .C(n538), .D(g1601), .Q(g6501)
         );
  AO22X1 U2752 ( .A(g1499), .B(n1167), .C(n539), .D(g1531), .Q(g6528)
         );
  AO22X1 U2753 ( .A(g1520), .B(n1169), .C(n538), .D(g1571), .Q(g6469)
         );
  AO22X1 U2754 ( .A(g1428), .B(n1169), .C(n538), .D(g1589), .Q(g6524)
         );
  AO22X1 U2755 ( .A(g1453), .B(n1167), .C(n539), .D(g1564), .Q(g6546)
         );
  AO22X1 U2756 ( .A(g1444), .B(n1169), .C(n538), .D(g1604), .Q(g6507)
         );
  AO22X1 U2757 ( .A(g1494), .B(n1167), .C(n539), .D(g1534), .Q(g6533)
         );
  AO22X1 U2758 ( .A(g1482), .B(n1167), .C(n539), .D(g1543), .Q(g6545)
         );
  AO22X1 U2759 ( .A(g1411), .B(n1169), .C(n538), .D(g1580), .Q(g6500)
         );
  AO22X1 U2760 ( .A(g1515), .B(n1169), .C(n538), .D(g1574), .Q(g6478)
         );
  AO22X1 U2761 ( .A(g1462), .B(n1167), .C(n539), .D(g1558), .Q(g6538)
         );
  AO22X1 U2762 ( .A(n624), .B(g1923), .C(n1039), .D(g1932), .Q(g8286)
         );
  AO22X1 U2763 ( .A(n650), .B(g709), .C(n1035), .D(g718), .Q(g8433) );
  AO22X1 U2764 ( .A(g166), .B(n1142), .C(n517), .D(g299), .Q(g6923) );
  AO22X1 U2765 ( .A(g178), .B(n1142), .C(n517), .D(g266), .Q(g6900) );
  AO22X1 U2766 ( .A(g158), .B(n1142), .C(n517), .D(g275), .Q(g6915) );
  AO22X1 U2767 ( .A(g182), .B(n1142), .C(n517), .D(g263), .Q(g6897) );
  AO22X1 U2768 ( .A(g153), .B(n1142), .C(n517), .D(g272), .Q(g6910) );
  AO22X1 U2769 ( .A(g139), .B(n1142), .C(n517), .D(g296), .Q(g6916) );
  AO22X1 U2770 ( .A(g127), .B(n1142), .C(n517), .D(g287), .Q(g6901) );
  AO22X1 U2771 ( .A(g131), .B(n1142), .C(n517), .D(g290), .Q(g6907) );
  AO22X1 U2772 ( .A(g143), .B(n1142), .C(n517), .D(g302), .Q(g6929) );
  AO22X1 U2773 ( .A(g135), .B(n1142), .C(n517), .D(g293), .Q(g6911) );
  AO22X1 U2774 ( .A(g148), .B(n1142), .C(n517), .D(g269), .Q(g6906) );
  AO22X1 U2775 ( .A(g174), .B(n1142), .C(n517), .D(g281), .Q(g6928) );
  AO22X1 U2776 ( .A(g170), .B(n1142), .C(n517), .D(g284), .Q(g6934) );
  AO22X1 U2777 ( .A(g162), .B(n1142), .C(n517), .D(g278), .Q(g6922) );
  AO22X1 U2778 ( .A(n954), .B(n1017), .C(n1018), .D(n668), .Q(g8631)
         );
  AO221X1 U2779 ( .A(n1027), .B(n1028), .C(n1029), .D(n1030), .E(
        n1716), .Q(n1017) );
  AO22X1 U2780 ( .A(n720), .B(n1713), .C(g636), .D(n1019), .Q(n1018)
         );
  AO22X1 U2781 ( .A(n624), .B(g1887), .C(n1039), .D(g1896), .Q(g8282)
         );
  AO22X1 U2782 ( .A(n650), .B(g673), .C(n1035), .D(g682), .Q(g8429) );
  AO22X1 U2783 ( .A(n650), .B(g718), .C(g727), .D(n1035), .Q(g8434) );
  AO22X1 U2784 ( .A(n624), .B(g1914), .C(n1039), .D(g1923), .Q(g8285)
         );
  AO22X1 U2785 ( .A(n624), .B(g1932), .C(g1941), .D(n1039), .Q(g8287)
         );
  AO22X1 U2786 ( .A(n650), .B(g700), .C(n1035), .D(g709), .Q(g8432) );
  AO22X1 U2787 ( .A(g351), .B(n1875), .C(g1083), .D(n1888), .Q(g6068)
         );
  AO22X1 U2788 ( .A(g336), .B(n1875), .C(test_so7), .D(n1888), .Q(
        g6054) );
  AO22X1 U2789 ( .A(g339), .B(n1875), .C(g1071), .D(n1888), .Q(g5910)
         );
  AO22X1 U2790 ( .A(g357), .B(n1875), .C(g1089), .D(n1888), .Q(g6080)
         );
  AO22X1 U2791 ( .A(g348), .B(n1875), .C(g1080), .D(n1888), .Q(g6059)
         );
  AO22X1 U2792 ( .A(g342), .B(n1875), .C(g1074), .D(n1888), .Q(g6099)
         );
  AO22X1 U2793 ( .A(g354), .B(n1875), .C(g1086), .D(n1888), .Q(g6071)
         );
  AO22X1 U2794 ( .A(g366), .B(n1875), .C(g1098), .D(n1888), .Q(g6096)
         );
  AO22X1 U2795 ( .A(g363), .B(n1875), .C(g1095), .D(n1888), .Q(g6093)
         );
  AO22X1 U2796 ( .A(g345), .B(n1875), .C(g1077), .D(n1888), .Q(g5914)
         );
  AO22X1 U2797 ( .A(g360), .B(n1875), .C(g1092), .D(n1888), .Q(g6088)
         );
  AO22X1 U2798 ( .A(g1621), .B(n1931), .C(n1955), .D(n986), .Q(g8771)
         );
  AO22X1 U2799 ( .A(g1630), .B(n1933), .C(n1955), .D(n971), .Q(g8776)
         );
  AO22X1 U2800 ( .A(g1615), .B(n1931), .C(n1955), .D(n987), .Q(g8770)
         );
  AO22X1 U2801 ( .A(g1512), .B(n1931), .C(n1955), .D(n1047), .Q(g8194)
         );
  XOR2X1 U2802 ( .A(n1596), .B(n1048), .Q(n1047) );
  NAND4X1 U2803 ( .A(g1104), .B(g1110), .C(n1654), .D(n1614), .Q(
        n1048) );
  AO22X1 U2804 ( .A(g1636), .B(n1924), .C(n1954), .D(n969), .Q(g8779)
         );
  AO22X1 U2805 ( .A(g1624), .B(n1932), .C(n1955), .D(n979), .Q(g8773)
         );
  AO22X1 U2806 ( .A(g1627), .B(n1932), .C(n1955), .D(n973), .Q(g8774)
         );
  AO22X1 U2807 ( .A(g1633), .B(n1931), .C(n1955), .D(n970), .Q(g8777)
         );
  AO22X1 U2808 ( .A(g4), .B(n1975), .C(n1161), .D(n1162), .Q(g6656) );
  NOR2X1 U2809 ( .A(n1163), .B(n1164), .Q(n1162) );
  NOR4X1 U2810 ( .A(n1165), .B(n1707), .C(n1166), .D(n1628), .Q(n1161) );
  OR4X1 U2811 ( .A(g1466), .B(g1482), .C(g1486), .D(g1499), .Q(n1163)
         );
  AO22X1 U2812 ( .A(n650), .B(g682), .C(n1035), .D(g691), .Q(g8430) );
  AO22X1 U2813 ( .A(n624), .B(g1896), .C(n1039), .D(g1905), .Q(g8283)
         );
  AO22X1 U2814 ( .A(n650), .B(g691), .C(n1035), .D(g700), .Q(g8431) );
  AO22X1 U2815 ( .A(n624), .B(g1905), .C(n1039), .D(g1914), .Q(g8284)
         );
  AO22X1 U2816 ( .A(n650), .B(g664), .C(n1035), .D(g673), .Q(g8428) );
  AO22X1 U2817 ( .A(n624), .B(g1878), .C(n1039), .D(g1887), .Q(g8281)
         );
  AO22X1 U2818 ( .A(test_so7), .B(n1954), .C(g1027), .D(n1934), .Q(
        g6894) );
  AO22X1 U2819 ( .A(g1710), .B(n1954), .C(g1713), .D(n1933), .Q(g5396)
         );
  AO22X1 U2820 ( .A(g1080), .B(n1953), .C(g995), .D(n1936), .Q(g6895)
         );
  AO22X1 U2821 ( .A(g1083), .B(n1953), .C(g991), .D(n1934), .Q(g6898)
         );
  AO22X1 U2822 ( .A(g1089), .B(n1953), .C(test_so8), .D(n1935), .Q(
        g6908) );
  AO22X1 U2823 ( .A(g1086), .B(n1953), .C(g1003), .D(n1935), .Q(g6902)
         );
  AO22X1 U2824 ( .A(g1077), .B(n1953), .C(g1032), .D(n1938), .Q(g7257)
         );
  AO22X1 U2825 ( .A(g1071), .B(n1953), .C(g1023), .D(n1939), .Q(g7244)
         );
  AO22X1 U2826 ( .A(g1092), .B(n1953), .C(g1011), .D(n1938), .Q(g6912)
         );
  AO22X1 U2827 ( .A(g1074), .B(n1953), .C(g1015), .D(n1939), .Q(g6930)
         );
  AO22X1 U2828 ( .A(n1885), .B(n1953), .C(g1718), .D(n1937), .Q(g5404)
         );
  AO22X1 U2829 ( .A(g1095), .B(n1953), .C(test_so2), .D(n1936), .Q(
        g6918) );
  AO22X1 U2830 ( .A(g1098), .B(n1953), .C(g1019), .D(n1937), .Q(g6924)
         );
  AO22X1 U2831 ( .A(g1941), .B(n624), .C(n1039), .D(g1950), .Q(g8288)
         );
  AO22X1 U2832 ( .A(g727), .B(n650), .C(n1035), .D(g736), .Q(g8435) );
  AO21X1 U2833 ( .A(g1615), .B(n1958), .C(n565), .Q(n1067) );
  AO21X1 U2834 ( .A(g1621), .B(n1958), .C(n564), .Q(n1075) );
  AO21X1 U2835 ( .A(g1624), .B(n1959), .C(n563), .Q(n1080) );
  AO21X1 U2836 ( .A(g1639), .B(n1959), .C(n566), .Q(n1063) );
  AO21X1 U2837 ( .A(g1618), .B(n1958), .C(n567), .Q(n1084) );
  NAND3X1 U2838 ( .A(g611), .B(n1645), .C(g591), .Q(n805) );
  AO21X1 U2839 ( .A(g566), .B(n1958), .C(n568), .Q(g6035) );
  AO21X1 U2840 ( .A(g554), .B(n1958), .C(n566), .Q(g6000) );
  AO21X1 U2841 ( .A(g560), .B(n1958), .C(n564), .Q(g6015) );
  AO21X1 U2842 ( .A(g546), .B(n1958), .C(n567), .Q(g5996) );
  AO21X1 U2843 ( .A(g557), .B(n1958), .C(n565), .Q(g6002) );
  AO21X1 U2844 ( .A(g569), .B(n1958), .C(n569), .Q(g6038) );
  AO21X1 U2845 ( .A(g563), .B(n1958), .C(n563), .Q(g6026) );
  ISOLANDX1 U2846 ( .D(g4175), .ISO(n1214), .Q(n1193) );
  ISOLANDX1 U2847 ( .D(g4177), .ISO(n1153), .Q(n1125) );
  ISOLANDX1 U2848 ( .D(g4179), .ISO(n1099), .Q(n1093) );
  AO221X1 U2849 ( .A(g1878), .B(n1031), .C(g1950), .D(n624), .E(
        n1032), .Q(g8559) );
  AO221X1 U2850 ( .A(g664), .B(n1016), .C(g736), .D(n650), .E(n954), 
        .Q(g8649) );
  AO221X1 U2851 ( .A(n1104), .B(n959), .C(g639), .D(n649), .E(n954), 
        .Q(g7626) );
  NOR2X1 U2852 ( .A(g639), .B(n1105), .Q(n1104) );
  NOR4X1 U2853 ( .A(n719), .B(n720), .C(n834), .D(n717), .Q(n1105) );
  NAND2X1 U2854 ( .A(g682), .B(n899), .Q(n957) );
  NAND2X1 U2855 ( .A(g1896), .B(n853), .Q(n896) );
  NAND2X1 U2856 ( .A(g1905), .B(n853), .Q(n890) );
  NAND2X1 U2857 ( .A(g691), .B(n899), .Q(n948) );
  NAND3X1 U2858 ( .A(g374), .B(g369), .C(g378), .Q(n1385) );
  ISOLANDX1 U2859 ( .D(n1137), .ISO(g12), .Q(n1159) );
  ISOLANDX1 U2860 ( .D(g810), .ISO(n1151), .Q(n1123) );
  ISOLANDX1 U2861 ( .D(g818), .ISO(n1097), .Q(n1090) );
  XOR3X1 U2862 ( .A(n1869), .B(g1003), .C(n1870), .Q(n1398) );
  XNOR2X1 U2863 ( .A(g1015), .B(g1011), .Q(n1870) );
  NAND2X1 U2864 ( .A(g1700), .B(DFF_275_n1), .Q(g4089) );
  XOR3X1 U2865 ( .A(n1871), .B(g1019), .C(n1872), .Q(n1397) );
  XNOR2X1 U2866 ( .A(test_so8), .B(g995), .Q(n1872) );
  ISOLANDX1 U2867 ( .D(n817), .ISO(g1834), .Q(n1380) );
  NAND2X1 U2868 ( .A(n555), .B(g1766), .Q(n1175) );
  NAND2X1 U2869 ( .A(n1191), .B(g806), .Q(n1151) );
  NAND2X1 U2870 ( .A(n1123), .B(g814), .Q(n1097) );
  NOR2X1 U2871 ( .A(n1873), .B(n711), .Q(g4904) );
  NOR2X1 U2872 ( .A(n1874), .B(n667), .Q(g4892) );
  AND2X1 U2873 ( .A(g1703), .B(n560), .Q(n1875) );
  NAND3X1 U2874 ( .A(n906), .B(n908), .C(g722), .Q(n902) );
  NAND3X1 U2875 ( .A(n861), .B(n863), .C(g1936), .Q(n857) );
  NAND3X1 U2876 ( .A(n718), .B(n1693), .C(n907), .Q(n901) );
  NAND3X1 U2877 ( .A(n712), .B(n1694), .C(n862), .Q(n856) );
  AND4X1 U2878 ( .A(g658), .B(n934), .C(g668), .D(n967), .Q(n906) );
  ISOLANDX1 U2879 ( .D(g713), .ISO(n1656), .Q(n967) );
  AND4X1 U2880 ( .A(g1872), .B(n876), .C(g1882), .D(n921), .Q(n861) );
  ISOLANDX1 U2881 ( .D(g1927), .ISO(n1657), .Q(n921) );
  ISOLANDX1 U2882 ( .D(g1160), .ISO(n1967), .Q(g4334) );
  ISOLANDX1 U2883 ( .D(g1166), .ISO(n1967), .Q(g4325) );
  ISOLANDX1 U2884 ( .D(g148), .ISO(n1967), .Q(g6759) );
  ISOLANDX1 U2885 ( .D(g1157), .ISO(n1967), .Q(g4338) );
  ISOLANDX1 U2886 ( .D(g1163), .ISO(n1967), .Q(g4330) );
  ISOLANDX1 U2887 ( .D(g237), .ISO(n1967), .Q(g6821) );
  ISOLANDX1 U2888 ( .D(g1499), .ISO(n1967), .Q(g6198) );
  ISOLANDX1 U2889 ( .D(g1411), .ISO(n1967), .Q(g6244) );
  ISOLANDX1 U2890 ( .D(g225), .ISO(n1967), .Q(g6826) );
  ISOLANDX1 U2891 ( .D(g1407), .ISO(n1967), .Q(g6216) );
  ISOLANDX1 U2892 ( .D(g213), .ISO(n1966), .Q(g6829) );
  ISOLANDX1 U2893 ( .D(g186), .ISO(n1966), .Q(g6833) );
  ISOLANDX1 U2894 ( .D(g219), .ISO(n1966), .Q(g6827) );
  ISOLANDX1 U2895 ( .D(g143), .ISO(n1966), .Q(g6757) );
  ISOLANDX1 U2896 ( .D(g207), .ISO(n1966), .Q(g6831) );
  ISOLANDX1 U2897 ( .D(g231), .ISO(n1966), .Q(g6822) );
  ISOLANDX1 U2898 ( .D(g192), .ISO(n1966), .Q(g6838) );
  ISOLANDX1 U2899 ( .D(test_so3), .ISO(n1966), .Q(g6823) );
  ISOLANDX1 U2900 ( .D(g1371), .ISO(n1966), .Q(g6824) );
  ISOLANDX1 U2901 ( .D(g1383), .ISO(n1966), .Q(g6832) );
  ISOLANDX1 U2902 ( .D(g243), .ISO(n1966), .Q(g6819) );
  NOR2X1 U2903 ( .A(g1878), .B(n622), .Q(n922) );
  NOR2X1 U2904 ( .A(g664), .B(n648), .Q(n846) );
  AO21X1 U2905 ( .A(g119), .B(n1969), .C(n1195), .Q(g5918) );
  AO21X1 U2906 ( .A(g12), .B(n1969), .C(n1195), .Q(g5445) );
  AO21X1 U2907 ( .A(g9), .B(n1974), .C(n1195), .Q(g5421) );
  AO21X1 U2908 ( .A(n597), .B(n884), .C(n596), .Q(g8939) );
  XNOR2X1 U2909 ( .A(g1909), .B(n885), .Q(n884) );
  NAND2X1 U2910 ( .A(n855), .B(n886), .Q(n885) );
  AO222X1 U2911 ( .A(n875), .B(g1900), .C(n877), .D(n1675), .E(g1914), .F(n853), .Q(n886) );
  AO21X1 U2912 ( .A(n605), .B(n897), .C(n606), .Q(g8926) );
  XOR2X1 U2913 ( .A(g731), .B(n898), .Q(n897) );
  OA221X1 U2914 ( .A(g736), .B(n648), .C(n899), .D(n900), .E(n850), 
        .Q(n898) );
  NAND2X1 U2915 ( .A(n901), .B(n902), .Q(n900) );
  AO21X1 U2916 ( .A(n605), .B(n903), .C(n606), .Q(g8923) );
  XOR2X1 U2917 ( .A(g722), .B(n904), .Q(n903) );
  OA221X1 U2918 ( .A(g727), .B(n648), .C(n905), .D(n899), .E(n850), 
        .Q(n904) );
  OA22X1 U2919 ( .A(n718), .B(n906), .C(n907), .D(n908), .Q(n905) );
  AO21X1 U2920 ( .A(n597), .B(n851), .C(n596), .Q(g8945) );
  XOR2X1 U2921 ( .A(g1945), .B(n852), .Q(n851) );
  OA221X1 U2922 ( .A(g1950), .B(n622), .C(n853), .D(n854), .E(n855), 
        .Q(n852) );
  NAND2X1 U2923 ( .A(n856), .B(n857), .Q(n854) );
  AO21X1 U2924 ( .A(n597), .B(n858), .C(n596), .Q(g8944) );
  XOR2X1 U2925 ( .A(g1936), .B(n859), .Q(n858) );
  OA221X1 U2926 ( .A(g1941), .B(n622), .C(n860), .D(n853), .E(n855), 
        .Q(n859) );
  OA22X1 U2927 ( .A(n712), .B(n861), .C(n862), .D(n863), .Q(n860) );
  AO21X1 U2928 ( .A(n597), .B(n872), .C(n596), .Q(g8941) );
  XNOR2X1 U2929 ( .A(g1927), .B(n873), .Q(n872) );
  NAND2X1 U2930 ( .A(n855), .B(n874), .Q(n873) );
  AO222X1 U2931 ( .A(n875), .B(n876), .C(n877), .D(n878), .E(g1932), 
        .F(n853), .Q(n874) );
  AO21X1 U2932 ( .A(n1182), .B(n1029), .C(n1042), .Q(g6243) );
  OR2X1 U2933 ( .A(g798), .B(g794), .Q(n1182) );
  OA22X1 U2934 ( .A(g639), .B(n1024), .C(n1692), .D(n1025), .Q(n1023)
         );
  NOR3X1 U2935 ( .A(n1655), .B(g1840), .C(n1608), .Q(n809) );
  OR4X1 U2936 ( .A(g1240), .B(g1245), .C(g1235), .D(n1330), .Q(n1329)
         );
  OR3X1 U2937 ( .A(g1250), .B(g1260), .C(g1255), .Q(n1330) );
  OR4X1 U2938 ( .A(g391), .B(g396), .C(g386), .D(n1438), .Q(n1437) );
  OR3X1 U2939 ( .A(g401), .B(g411), .C(g406), .Q(n1438) );
  NAND2X1 U2940 ( .A(n1969), .B(n1058), .Q(n1040) );
  NAND3X1 U2941 ( .A(DFF_436_n1), .B(n594), .C(n1059), .Q(n1058) );
  NAND2X1 U2942 ( .A(n1969), .B(n1235), .Q(n1224) );
  NAND3X1 U2943 ( .A(n1236), .B(n1683), .C(g1212), .Q(n1235) );
  NAND2X1 U2944 ( .A(n1090), .B(g822), .Q(n1043) );
  NBUFFX1 U2945 ( .IN(g1713), .Q(n1885) );
  NAND2X1 U2946 ( .A(n520), .B(g794), .Q(g5849) );
  NAND3X1 U2947 ( .A(n804), .B(g605), .C(n721), .Q(n837) );
  AOI22X1 U2948 ( .A(n1876), .B(n1877), .C(n1878), .D(g431), .Q(n1434) );
  OAI21X1 U2949 ( .A(n1436), .B(n1437), .C(n1878), .Q(n1877) );
  OA21X1 U2950 ( .A(n1052), .B(n1053), .C(n1610), .Q(g8173) );
  OA21X1 U2951 ( .A(n1054), .B(n1055), .C(g1806), .Q(n1053) );
  AND3X1 U2952 ( .A(n1056), .B(n1055), .C(g1801), .Q(n1052) );
  NAND3X1 U2953 ( .A(g1801), .B(n1057), .C(g1806), .Q(n1055) );
  OR4X1 U2954 ( .A(test_so6), .B(g1275), .C(g1265), .D(n1331), .Q(
        n1328) );
  OR4X1 U2955 ( .A(g1304), .B(g1300), .C(g1296), .D(g1292), .Q(n1331)
         );
  OR4X1 U2956 ( .A(g421), .B(g426), .C(g416), .D(n1439), .Q(n1436) );
  OR4X1 U2957 ( .A(g452), .B(g448), .C(g444), .D(g440), .Q(n1439) );
  NOR2X1 U2958 ( .A(n1041), .B(n1042), .Q(g8245) );
  XOR2X1 U2959 ( .A(n1043), .B(g826), .Q(n1041) );
  OAI22X1 U2960 ( .A(g525), .B(n1698), .C(g521), .D(n1354), .Q(n1241)
         );
  OA21X1 U2961 ( .A(n1355), .B(n1356), .C(n1695), .Q(n1354) );
  NOR2X1 U2962 ( .A(n954), .B(n961), .Q(g8820) );
  XOR2X1 U2963 ( .A(n603), .B(g622), .Q(n961) );
  NAND3X1 U2964 ( .A(g4892), .B(n1020), .C(n1021), .Q(n1019) );
  NAND4X1 U2965 ( .A(n1024), .B(n1026), .C(n953), .D(n1025), .Q(n1020) );
  XOR2X1 U2966 ( .A(n1022), .B(n1023), .Q(n1021) );
  NAND2X1 U2967 ( .A(g255), .B(g622), .Q(n1022) );
  NAND3X1 U2968 ( .A(n1118), .B(n1119), .C(n643), .Q(g7441) );
  NAND2X1 U2969 ( .A(g643), .B(n1701), .Q(n1118) );
  INVX1 U2970 ( .IN(n1101), .Q(n643) );
  NOR2X1 U2971 ( .A(n1964), .B(n1062), .Q(g8055) );
  XNOR2X1 U2972 ( .A(g1490), .B(n1063), .Q(n1062) );
  NOR2X1 U2973 ( .A(n1963), .B(n1078), .Q(g8044) );
  XNOR2X1 U2974 ( .A(g131), .B(g6038), .Q(n1078) );
  NOR2X1 U2975 ( .A(n1964), .B(n1064), .Q(g8054) );
  XNOR2X1 U2976 ( .A(g174), .B(g6015), .Q(n1064) );
  NOR2X1 U2977 ( .A(n1983), .B(n1065), .Q(g8053) );
  XNOR2X1 U2978 ( .A(g139), .B(g6045), .Q(n1065) );
  NOR2X1 U2979 ( .A(n1964), .B(n1061), .Q(g8059) );
  XNOR2X1 U2980 ( .A(g135), .B(g6042), .Q(n1061) );
  NOR2X1 U2981 ( .A(n1983), .B(n1066), .Q(g8052) );
  XNOR2X1 U2982 ( .A(g1486), .B(n1067), .Q(n1066) );
  NOR2X1 U2983 ( .A(n1966), .B(n1071), .Q(g8049) );
  XNOR2X1 U2984 ( .A(g166), .B(g6049), .Q(n1071) );
  NOR2X1 U2985 ( .A(n1983), .B(n1072), .Q(g8048) );
  XNOR2X1 U2986 ( .A(g153), .B(g5996), .Q(n1072) );
  NOR2X1 U2987 ( .A(n1962), .B(n1079), .Q(g8043) );
  XNOR2X1 U2988 ( .A(g1478), .B(n1080), .Q(n1079) );
  NOR2X1 U2989 ( .A(n1962), .B(n1085), .Q(g8040) );
  XNOR2X1 U2990 ( .A(g1474), .B(n1086), .Q(n1085) );
  NOR2X1 U2991 ( .A(n1963), .B(n972), .Q(g8775) );
  XNOR2X1 U2992 ( .A(g1436), .B(n973), .Q(n972) );
  NOR2X1 U2993 ( .A(n1964), .B(n1060), .Q(g8060) );
  XNOR2X1 U2994 ( .A(g162), .B(g6002), .Q(n1060) );
  NOR2X1 U2995 ( .A(n1962), .B(n1087), .Q(g8039) );
  XNOR2X1 U2996 ( .A(g1470), .B(n1088), .Q(n1087) );
  NOR2X1 U2997 ( .A(n1962), .B(n1095), .Q(g7843) );
  XNOR2X1 U2998 ( .A(g158), .B(g6000), .Q(n1095) );
  NOR2X1 U2999 ( .A(n1962), .B(n1076), .Q(g8045) );
  XNOR2X1 U3000 ( .A(g1462), .B(n1077), .Q(n1076) );
  NOR2X1 U3001 ( .A(n1962), .B(n988), .Q(g8769) );
  XNOR2X1 U3002 ( .A(g1428), .B(n987), .Q(n988) );
  NOR2X1 U3003 ( .A(n1983), .B(n1070), .Q(g8050) );
  XNOR2X1 U3004 ( .A(g170), .B(g6026), .Q(n1070) );
  NOR2X1 U3005 ( .A(n1983), .B(n1068), .Q(g8051) );
  XNOR2X1 U3006 ( .A(g1466), .B(n1069), .Q(n1068) );
  NOR2X1 U3007 ( .A(n1962), .B(n1074), .Q(g8046) );
  XNOR2X1 U3008 ( .A(g1482), .B(n1075), .Q(n1074) );
  NOR2X1 U3009 ( .A(n1966), .B(n1006), .Q(g8766) );
  XNOR2X1 U3010 ( .A(g1448), .B(n969), .Q(n1006) );
  NOR2X1 U3011 ( .A(n1962), .B(n1083), .Q(g8041) );
  XNOR2X1 U3012 ( .A(g1494), .B(n1084), .Q(n1083) );
  NBUFFX1 U3013 ( .IN(g1690), .Q(n1882) );
  NOR2X1 U3014 ( .A(n1961), .B(n994), .Q(g8768) );
  XNOR2X1 U3015 ( .A(g1444), .B(n970), .Q(n994) );
  NOR2X1 U3016 ( .A(n1961), .B(n1011), .Q(g8765) );
  XNOR2X1 U3017 ( .A(g1432), .B(n979), .Q(n1011) );
  NOR2X1 U3018 ( .A(n1961), .B(n1000), .Q(g8767) );
  XNOR2X1 U3019 ( .A(g1403), .B(n986), .Q(n1000) );
  NOR2X1 U3020 ( .A(n1961), .B(n980), .Q(g8772) );
  XNOR2X1 U3021 ( .A(g1440), .B(n971), .Q(n980) );
  NOR4X1 U3022 ( .A(n1275), .B(n1276), .C(n1277), .D(n1278), .Q(n1274) );
  XOR2X1 U3023 ( .A(test_so8), .B(g1245), .Q(n1276) );
  XOR2X1 U3024 ( .A(g991), .B(g1235), .Q(n1278) );
  XOR2X1 U3025 ( .A(g1250), .B(g1011), .Q(n1277) );
  NOR4X1 U3026 ( .A(n1425), .B(n1426), .C(n1427), .D(n1428), .Q(n1424) );
  XOR2X1 U3027 ( .A(g396), .B(g324), .Q(n1426) );
  XOR2X1 U3028 ( .A(g386), .B(g318), .Q(n1428) );
  XOR2X1 U3029 ( .A(g401), .B(g327), .Q(n1427) );
  NOR4X1 U3030 ( .A(g1166), .B(g1163), .C(g1160), .D(g1157), .Q(n1269) );
  NBUFFX1 U3031 ( .IN(g456), .Q(n1884) );
  NOR3X1 U3032 ( .A(g1909), .B(g1918), .C(g1900), .Q(n878) );
  NOR3X1 U3033 ( .A(g695), .B(g704), .C(g686), .Q(n936) );
  NOR3X1 U3034 ( .A(g1861), .B(g1864), .C(n1642), .Q(n1147) );
  NOR2X1 U3035 ( .A(n711), .B(DFF_489_n1), .Q(g4905) );
  NOR2X1 U3036 ( .A(n711), .B(DFF_385_n1), .Q(g4902) );
  NOR2X1 U3037 ( .A(n711), .B(DFF_330_n1), .Q(g4903) );
  NOR2X1 U3038 ( .A(n667), .B(DFF_157_n1), .Q(g4893) );
  NOR2X1 U3039 ( .A(n667), .B(DFF_336_n1), .Q(g4890) );
  NOR2X1 U3040 ( .A(n667), .B(DFF_136_n1), .Q(g4891) );
  NOR2X1 U3041 ( .A(n1199), .B(n1961), .Q(g5755) );
  XOR3X1 U3042 ( .A(g1389), .B(n1200), .C(n1201), .Q(n1199) );
  XOR2X1 U3043 ( .A(g201), .B(g197), .Q(n1201) );
  NOR2X1 U3044 ( .A(g1386), .B(n1202), .Q(n1200) );
  NOR2X1 U3045 ( .A(n1179), .B(n1961), .Q(g6439) );
  XNOR3X1 U3046 ( .A(n1180), .B(g153), .C(g182), .Q(n1179) );
  XOR2X1 U3047 ( .A(g148), .B(g143), .Q(n1180) );
  NOR2X1 U3048 ( .A(n1196), .B(n1961), .Q(g5770) );
  XOR3X1 U3049 ( .A(n1197), .B(g1499), .C(n1707), .Q(n1196) );
  XOR2X1 U3050 ( .A(g1494), .B(g1453), .Q(n1197) );
  OR2X1 U3051 ( .A(g1900), .B(g1909), .Q(n882) );
  OR2X1 U3052 ( .A(g686), .B(g695), .Q(n940) );
  NAND2X1 U3053 ( .A(n995), .B(n996), .Q(n970) );
  AO221X1 U3054 ( .A(n997), .B(g1141), .C(n1660), .D(n998), .E(g2355), .Q(n996) );
  NOR2X1 U3055 ( .A(g1101), .B(n999), .Q(n997) );
  NAND2X1 U3056 ( .A(n634), .B(n1654), .Q(n998) );
  NAND2X1 U3057 ( .A(n981), .B(n982), .Q(n971) );
  AO221X1 U3058 ( .A(n983), .B(g1137), .C(n1597), .D(n984), .E(g2355), .Q(n982) );
  NAND2X1 U3059 ( .A(n631), .B(g1101), .Q(n984) );
  NOR2X1 U3060 ( .A(n1654), .B(n978), .Q(n983) );
  NAND2X1 U3061 ( .A(n989), .B(n990), .Q(n987) );
  AO221X1 U3062 ( .A(n991), .B(g1121), .C(n1618), .D(n992), .E(g2355), .Q(n990) );
  NOR2X1 U3063 ( .A(n1654), .B(n993), .Q(n991) );
  NAND2X1 U3064 ( .A(n632), .B(g1101), .Q(n992) );
  AND4X1 U3065 ( .A(n1625), .B(n1688), .C(n1208), .D(n1209), .Q(n1184)
         );
  NOR2X1 U3066 ( .A(g1371), .B(test_so3), .Q(n1208) );
  NOR4X1 U3067 ( .A(g243), .B(g237), .C(g231), .D(g225), .Q(n1209) );
  AO21X1 U3068 ( .A(n605), .B(n942), .C(n606), .Q(g8887) );
  XNOR2X1 U3069 ( .A(g695), .B(n943), .Q(n942) );
  NAND2X1 U3070 ( .A(n850), .B(n944), .Q(n943) );
  AO222X1 U3071 ( .A(n933), .B(g686), .C(n935), .D(n1676), .E(g700), 
        .F(n899), .Q(n944) );
  NOR2X1 U3072 ( .A(n1191), .B(n1212), .Q(g5543) );
  OA22X1 U3073 ( .A(n1622), .B(n1042), .C(g5849), .D(n1717), .Q(n1212)
         );
  XNOR2X1 U3074 ( .A(test_so1), .B(n1045), .Q(N599) );
  NOR3X1 U3075 ( .A(g1125), .B(g1133), .C(g1129), .Q(n1268) );
  AO21X1 U3076 ( .A(n597), .B(n879), .C(n596), .Q(g8940) );
  XOR2X1 U3077 ( .A(g1918), .B(n880), .Q(n879) );
  NOR2X1 U3078 ( .A(n881), .B(n620), .Q(n880) );
  OA222X1 U3079 ( .A(n622), .B(n1718), .C(n600), .D(n882), .E(n595), 
        .F(n883), .Q(n881) );
  AO21X1 U3080 ( .A(n605), .B(n937), .C(n606), .Q(g8889) );
  XOR2X1 U3081 ( .A(g704), .B(n938), .Q(n937) );
  NOR2X1 U3082 ( .A(n939), .B(n644), .Q(n938) );
  OA222X1 U3083 ( .A(n648), .B(n1719), .C(n645), .D(n940), .E(n646), 
        .F(n941), .Q(n939) );
  NOR3X1 U3084 ( .A(n1431), .B(n1432), .C(n1433), .Q(n1423) );
  XOR2X1 U3085 ( .A(g421), .B(g312), .Q(n1431) );
  XOR2X1 U3086 ( .A(g411), .B(g333), .Q(n1433) );
  XOR2X1 U3087 ( .A(n1681), .B(n1390), .Q(n1432) );
  NBUFFX1 U3088 ( .IN(g456), .Q(n1883) );
  NOR3X1 U3089 ( .A(n1150), .B(n1123), .C(n1042), .Q(g6733) );
  ISOLANDX1 U3090 ( .D(n1151), .ISO(g810), .Q(n1150) );
  NOR3X1 U3091 ( .A(n1096), .B(n1090), .C(n1042), .Q(g7709) );
  ISOLANDX1 U3092 ( .D(n1097), .ISO(g818), .Q(n1096) );
  NOR3X1 U3093 ( .A(n1098), .B(n1093), .C(n537), .Q(g7705) );
  ISOLANDX1 U3094 ( .D(n1099), .ISO(g4179), .Q(n1098) );
  NOR3X1 U3095 ( .A(n1213), .B(n1193), .C(n537), .Q(g5536) );
  ISOLANDX1 U3096 ( .D(n1214), .ISO(g4175), .Q(n1213) );
  NOR3X1 U3097 ( .A(n1152), .B(n1125), .C(n537), .Q(g6728) );
  ISOLANDX1 U3098 ( .D(n1153), .ISO(g4177), .Q(n1152) );
  NAND4X1 U3099 ( .A(n1159), .B(g1470), .C(g1474), .D(g1494), .Q(
        n1165) );
  NBUFFX1 U3100 ( .IN(g1690), .Q(n1881) );
  NOR2X1 U3101 ( .A(n1885), .B(n1174), .Q(g6508) );
  OA22X1 U3102 ( .A(n1175), .B(n1176), .C(n553), .D(n1715), .Q(n1174)
         );
  NAND2X1 U3103 ( .A(test_so5), .B(n1172), .Q(n1176) );
  NOR2X1 U3104 ( .A(n1885), .B(n1138), .Q(g6983) );
  OA22X1 U3105 ( .A(n1139), .B(n1140), .C(n1116), .D(n1702), .Q(n1138)
         );
  NAND2X1 U3106 ( .A(g1786), .B(n1117), .Q(n1140) );
  NAND4X1 U3107 ( .A(n1679), .B(n1620), .C(n1600), .D(n1358), .Q(
        n1355) );
  NOR4X1 U3108 ( .A(g542), .B(g538), .C(g534), .D(g530), .Q(n1358) );
  NOR2X1 U3109 ( .A(n1885), .B(n1094), .Q(g7930) );
  XNOR2X1 U3110 ( .A(n1056), .B(g1801), .Q(n1094) );
  NOR2X1 U3111 ( .A(n1957), .B(n818), .Q(g9269) );
  XOR2X1 U3112 ( .A(g1822), .B(n819), .Q(n818) );
  NOR2X1 U3113 ( .A(n820), .B(n821), .Q(n819) );
  AOI21X1 U3114 ( .A(n822), .B(n815), .C(n598), .Q(n821) );
  NOR2X1 U3115 ( .A(n1958), .B(n1033), .Q(g8505) );
  XOR2X1 U3116 ( .A(g617), .B(n1034), .Q(n1033) );
  AOI21X1 U3117 ( .A(n650), .B(g736), .C(n960), .Q(n1034) );
  NOR2X1 U3118 ( .A(n1958), .B(n800), .Q(g9721) );
  XOR2X1 U3119 ( .A(g611), .B(n801), .Q(n800) );
  OA21X1 U3120 ( .A(n802), .B(n649), .C(n803), .Q(n801) );
  OA21X1 U3121 ( .A(n804), .B(n805), .C(n1645), .Q(n802) );
  NOR2X1 U3122 ( .A(n1957), .B(n835), .Q(g9124) );
  XOR2X1 U3123 ( .A(g599), .B(n836), .Q(n835) );
  ISOLANDX1 U3124 ( .D(n837), .ISO(n838), .Q(n836) );
  OA21X1 U3125 ( .A(n720), .B(n717), .C(n804), .Q(n838) );
  NOR2X1 U3126 ( .A(n1957), .B(n823), .Q(g9266) );
  XOR2X1 U3127 ( .A(g1814), .B(n824), .Q(n823) );
  NOR2X1 U3128 ( .A(n825), .B(n820), .Q(n824) );
  OA21X1 U3129 ( .A(n809), .B(n713), .C(n812), .Q(n825) );
  NOR2X1 U3130 ( .A(n1885), .B(n1177), .Q(g6502) );
  XOR2X1 U3131 ( .A(n1175), .B(test_so5), .Q(n1177) );
  NOR2X1 U3132 ( .A(n1885), .B(n1168), .Q(g6525) );
  XOR2X1 U3133 ( .A(n1139), .B(g1786), .Q(n1168) );
  NOR2X1 U3134 ( .A(n1958), .B(n1036), .Q(g8384) );
  XOR2X1 U3135 ( .A(g1840), .B(n1037), .Q(n1036) );
  AOI21X1 U3136 ( .A(n624), .B(g1950), .C(n929), .Q(n1037) );
  NAND4X1 U3137 ( .A(n1680), .B(n1621), .C(n1599), .D(n1357), .Q(
        n1356) );
  NOR3X1 U3138 ( .A(g491), .B(g501), .C(g496), .Q(n1357) );
  INVX1 U3139 ( .IN(g23), .Q(g3327) );
  INVX1 U3140 ( .IN(g18), .Q(n1960) );
  NAND2X1 U3141 ( .A(n1279), .B(n1280), .Q(n1275) );
  XNOR2X1 U3142 ( .A(g995), .B(g1275), .Q(n1279) );
  XNOR2X1 U3143 ( .A(g1003), .B(g1240), .Q(n1280) );
  NAND2X1 U3144 ( .A(n1429), .B(n1430), .Q(n1425) );
  XNOR2X1 U3145 ( .A(g315), .B(g426), .Q(n1429) );
  XNOR2X1 U3146 ( .A(g321), .B(g391), .Q(n1430) );
  INVX1 U3147 ( .IN(g881), .Q(n594) );
  NAND2X1 U3148 ( .A(g1703), .B(n1724), .Q(n1451) );
  NAND2X1 U3149 ( .A(n1229), .B(g1351), .Q(n1228) );
  NAND2X1 U3150 ( .A(n617), .B(g986), .Q(n1338) );
  AND3X1 U3151 ( .A(g1336), .B(g1346), .C(g1341), .Q(n1229) );
  NAND3X1 U3152 ( .A(n1612), .B(n1595), .C(g650), .Q(n1129) );
  NAND3X1 U3153 ( .A(g971), .B(g981), .C(g976), .Q(n1342) );
  NAND2X1 U3154 ( .A(g1909), .B(g1900), .Q(n883) );
  NAND2X1 U3155 ( .A(g695), .B(g686), .Q(n941) );
  AO22X1 U3156 ( .A(g1786), .B(n725), .C(g1750), .D(n1217), .Q(g4264)
         );
  AO22X1 U3157 ( .A(g1796), .B(n725), .C(g1756), .D(n1217), .Q(g4283)
         );
  AO22X1 U3158 ( .A(g1781), .B(n725), .C(g1747), .D(n1217), .Q(g4255)
         );
  AO22X1 U3159 ( .A(g1806), .B(n725), .C(g1762), .D(n1217), .Q(g4309)
         );
  AO22X1 U3160 ( .A(g1766), .B(n725), .C(g1738), .D(n1217), .Q(g4231)
         );
  AO22X1 U3161 ( .A(g1791), .B(n725), .C(g1753), .D(n1217), .Q(g4274)
         );
  AO22X1 U3162 ( .A(test_so5), .B(n725), .C(g1741), .D(n1217), .Q(
        g4238) );
  AO22X1 U3163 ( .A(g1801), .B(n725), .C(g1759), .D(n1217), .Q(g4293)
         );
  AO22X1 U3164 ( .A(g1776), .B(n725), .C(g1744), .D(n1217), .Q(g4239)
         );
  NAND4X1 U3165 ( .A(g1444), .B(g1428), .C(g1440), .D(g1436), .Q(
        n1157) );
  NAND4X1 U3166 ( .A(g1478), .B(g1462), .C(g1490), .D(n1703), .Q(
        n1164) );
  NAND2X1 U3167 ( .A(g806), .B(g802), .Q(n1030) );
  NOR2X1 U3168 ( .A(g1737), .B(g1610), .Q(g2478) );
  NOR2X1 U3169 ( .A(n562), .B(n1189), .Q(g6155) );
  XOR2X1 U3170 ( .A(g1707), .B(n1653), .Q(n1189) );
  ISOLANDX1 U3171 ( .D(g1610), .ISO(n555), .Q(g5194) );
  NAND2X1 U3172 ( .A(n1131), .B(n1610), .Q(g7133) );
  XOR2X1 U3173 ( .A(g1766), .B(n1054), .Q(n1131) );
  AO21X1 U3174 ( .A(g654), .B(n1100), .C(n1101), .Q(g7660) );
  NAND4X1 U3175 ( .A(g627), .B(n1612), .C(n1595), .D(n1709), .Q(n1100) );
  AO21X1 U3176 ( .A(g1868), .B(n1143), .C(n1144), .Q(g6909) );
  OR3X1 U3177 ( .A(g1861), .B(g1864), .C(n1642), .Q(n1143) );
  OA21X1 U3178 ( .A(n1146), .B(n1147), .C(n619), .Q(g6795) );
  OA21X1 U3179 ( .A(g1861), .B(n1642), .C(g1864), .Q(n1146) );
  OA21X1 U3180 ( .A(n1218), .B(n592), .C(g746), .Q(g3462) );
  NOR2X1 U3181 ( .A(g750), .B(n1647), .Q(n1218) );
  NOR2X1 U3182 ( .A(n1178), .B(n1144), .Q(g6471) );
  XOR2X1 U3183 ( .A(n1642), .B(g1861), .Q(n1178) );
  NOR4X1 U3184 ( .A(n1210), .B(n1211), .C(n1702), .D(n1626), .Q(g5556) );
  NAND4X1 U3185 ( .A(n1882), .B(g1707), .C(g1806), .D(g1801), .Q(
        n1210) );
  NAND3X1 U3186 ( .A(n661), .B(n1659), .C(g1786), .Q(n1211) );
  NOR2X1 U3187 ( .A(g1707), .B(n562), .Q(g4076) );
  NAND2X1 U3188 ( .A(g814), .B(g810), .Q(n1028) );
  NAND2X1 U3189 ( .A(g822), .B(g818), .Q(n1027) );
  NAND4X1 U3190 ( .A(g170), .B(g174), .C(n1613), .D(n1704), .Q(n1135)
         );
  OR2X1 U3191 ( .A(g1289), .B(g1212), .Q(g4556) );
  INVX1 U3192 ( .IN(g1700), .Q(n562) );
  AND2X1 U3193 (.A(g6179), .B(n519), .Q(Tg1_OUT1));
  AND2X1 U3194 (.A(n1202), .B(n1132), .Q(Tg1_OUT2));
  AND2X1 U3195 (.A(n1226), .B(n1858), .Q(Tg1_OUT3));
  AND2X1 U3196 (.A(g5556), .B(n898), .Q(Tg1_OUT4));
  AND4X1 U3197 (.A(Tg1_OUT1), .B(Tg1_OUT2), .C(Tg1_OUT3), .D(Tg1_OUT4), .Q(Tg1_OUT1234));
  NOR2X1 U3198 (.A(n1391), .B(n931), .Q(Tg1_OUT5));
  NOR2X1 U3199 (.A(n857), .B(n902), .Q(Tg1_OUT6));
  NOR2X1 U3200 (.A(n1889), .B(n1890), .Q(Tg1_OUT7));
  NOR2X1 U3201 (.A(n1055), .B(n1016), .Q(Tg1_OUT8));
  AND4X1 U3202 (.A(Tg1_OUT5), .B(Tg1_OUT6), .C(Tg1_OUT7), .D(Tg1_OUT8), .Q(Tg1_OUT5678));
  AND2X1 U3203 ( .A(Tg1_OUT1234), .B(Tg1_OUT5678), .Q(Tg1_Trigger1) );
  DFFNX2 U3204 ( .CLK(Tg1_Trigger1), .D(1'b1), .Q(Tg1) ); 
  AND2X1 U3205 (.A(n938), .B(n1917), .Q(Tg2_OUT1));
  AND2X1 U3206 (.A(n1921), .B(n1911), .Q(Tg2_OUT2));
  AND2X1 U3207 (.A(n1918), .B(n1913), .Q(Tg2_OUT3));
  AND2X1 U3208 (.A(n1916), .B(n1910), .Q(Tg2_OUT4));
  AND4X1 U3209 (.A(Tg2_OUT1), .B(Tg2_OUT2), .C(Tg2_OUT3), .D(Tg2_OUT4), .Q(Tg2_OUT1234));
  AND2X1 U3210 (.A(n1161), .B(n1154), .Q(Tg2_OUT5));
  AND2X1 U3211 (.A(n1116), .B(n1162), .Q(Tg2_OUT6));
  AND2X1 U3212 (.A(n1155), .B(n1107), .Q(Tg2_OUT7));
  AND2X1 U3213 (.A(n929), .B(n554), .Q(Tg2_OUT8));
  AND4X1 U3214 (.A(Tg2_OUT5), .B(Tg2_OUT6), .C(Tg2_OUT7), .D(Tg2_OUT8), .Q(Tg2_OUT5678));
  AND2X1 U3215 ( .A(Tg2_OUT1234), .B(Tg2_OUT5678), .Q(Tg2_Trigger2) );
  DFFNX2 U3216 ( .CLK(Tg2_Trigger2), .D(Tg1), .Q(Tg2) ); 
  INVX1 U3217 ( .IN(test_se), .Q(test_se_NOT) );
  AND2X1 U3218 (.A(Tg2), .B(test_se_NOT), .Q(Trigger_select) );
  MUX21X2 U3219 ( .A(g4207_Payload), .B(n1936), .S(Trigger_select), .Q(g4207) );

endmodule

