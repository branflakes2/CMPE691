library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity vigenere_encoder is

port
